----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 10/08/2020 06:37:32 PM
-- Design Name: 
-- Module Name: FIR_Example - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity FIR_Example is
	Generic(
		cIWGlobal		: integer := 32; --Input Integer part Width
		cFWGlobal		: integer := 32 --Input Fractional part Width
		);
    Port (
		--General Ports
		   Clk		: in STD_LOGIC;
		   Rst		: in STD_LOGIC;
		   
		--Functional Inputs
		--Input of the FIR Filter
		   X		: in Signed (cIWGlobal+cFWGlobal-1 downto 0);
		-- The Output of the FIR Filter
           Y		: out Signed (cIWGlobal+cFWGlobal-1 downto 0);
		
		
		--Width inputs
		   Add000aIW	: in integer range 0 to cIWGlobal;
		   Add001aIW	: in integer range 0 to cIWGlobal;
		   Add002aIW	: in integer range 0 to cIWGlobal;
		   Add003aIW	: in integer range 0 to cIWGlobal;
		   Add004aIW	: in integer range 0 to cIWGlobal;
		   Add005aIW	: in integer range 0 to cIWGlobal;
		   Add006aIW	: in integer range 0 to cIWGlobal;
		   Add007aIW	: in integer range 0 to cIWGlobal;
		   Add008aIW	: in integer range 0 to cIWGlobal;
		   Add009aIW	: in integer range 0 to cIWGlobal;
		   Add010aIW	: in integer range 0 to cIWGlobal;
		   Add011aIW	: in integer range 0 to cIWGlobal;
		   Add012aIW	: in integer range 0 to cIWGlobal;
		   Add013aIW	: in integer range 0 to cIWGlobal;
		   Add014aIW	: in integer range 0 to cIWGlobal;
		   Add015aIW	: in integer range 0 to cIWGlobal;
		   Add016aIW	: in integer range 0 to cIWGlobal;
		   Add017aIW	: in integer range 0 to cIWGlobal;
		   Add018aIW	: in integer range 0 to cIWGlobal;
		   Add019aIW	: in integer range 0 to cIWGlobal;
		   Add020aIW	: in integer range 0 to cIWGlobal;
		   Add021aIW	: in integer range 0 to cIWGlobal;
		   Add022aIW	: in integer range 0 to cIWGlobal;
		   Add023aIW	: in integer range 0 to cIWGlobal;
		   Add024aIW	: in integer range 0 to cIWGlobal;
		   Add025aIW	: in integer range 0 to cIWGlobal;
		   Add026aIW	: in integer range 0 to cIWGlobal;
		   Add027aIW	: in integer range 0 to cIWGlobal;
		   Add028aIW	: in integer range 0 to cIWGlobal;
		   Add029aIW	: in integer range 0 to cIWGlobal;
		   Add030aIW	: in integer range 0 to cIWGlobal;
		   Add031aIW	: in integer range 0 to cIWGlobal;
		   Add032aIW	: in integer range 0 to cIWGlobal;
		   Add033aIW	: in integer range 0 to cIWGlobal;
		   Add034aIW	: in integer range 0 to cIWGlobal;
		   Add035aIW	: in integer range 0 to cIWGlobal;
		   Add036aIW	: in integer range 0 to cIWGlobal;
		   Add037aIW	: in integer range 0 to cIWGlobal;
		   Add038aIW	: in integer range 0 to cIWGlobal;
		   Add039aIW	: in integer range 0 to cIWGlobal;
		   Add040aIW	: in integer range 0 to cIWGlobal;
		   Add041aIW	: in integer range 0 to cIWGlobal;
		   Add042aIW	: in integer range 0 to cIWGlobal;
		   Add043aIW	: in integer range 0 to cIWGlobal;
		   Add044aIW	: in integer range 0 to cIWGlobal;
		   Add045aIW	: in integer range 0 to cIWGlobal;
		   Add046aIW	: in integer range 0 to cIWGlobal;
		   Add047aIW	: in integer range 0 to cIWGlobal;
		   Add048aIW	: in integer range 0 to cIWGlobal;
		   Add049aIW	: in integer range 0 to cIWGlobal;
		   Add050aIW	: in integer range 0 to cIWGlobal;
		   Add051aIW	: in integer range 0 to cIWGlobal;
		   Add052aIW	: in integer range 0 to cIWGlobal;
		   Add053aIW	: in integer range 0 to cIWGlobal;
		   Add054aIW	: in integer range 0 to cIWGlobal;
		   Add055aIW	: in integer range 0 to cIWGlobal;
		   Add056aIW	: in integer range 0 to cIWGlobal;
		   Add057aIW	: in integer range 0 to cIWGlobal;
		   Add058aIW	: in integer range 0 to cIWGlobal;
		   Add059aIW	: in integer range 0 to cIWGlobal;
		   Add060aIW	: in integer range 0 to cIWGlobal;
		   Add061aIW	: in integer range 0 to cIWGlobal;
		   Add062aIW	: in integer range 0 to cIWGlobal;
		   Add063aIW	: in integer range 0 to cIWGlobal;
		   Add064aIW	: in integer range 0 to cIWGlobal;
		   Add065aIW	: in integer range 0 to cIWGlobal;
		   Add066aIW	: in integer range 0 to cIWGlobal;
		   Add067aIW	: in integer range 0 to cIWGlobal;
		   Add068aIW	: in integer range 0 to cIWGlobal;
		   Add069aIW	: in integer range 0 to cIWGlobal;
		   Add070aIW	: in integer range 0 to cIWGlobal;
		   Add071aIW	: in integer range 0 to cIWGlobal;
		   Add072aIW	: in integer range 0 to cIWGlobal;
		   Add073aIW	: in integer range 0 to cIWGlobal;
		   Add074aIW	: in integer range 0 to cIWGlobal;
		   Add075aIW	: in integer range 0 to cIWGlobal;
		   Add076aIW	: in integer range 0 to cIWGlobal;
		   Add077aIW	: in integer range 0 to cIWGlobal;
		   Add078aIW	: in integer range 0 to cIWGlobal;
		   Add079aIW	: in integer range 0 to cIWGlobal;
		   Add080aIW	: in integer range 0 to cIWGlobal;
		   Add081aIW	: in integer range 0 to cIWGlobal;
		   Add082aIW	: in integer range 0 to cIWGlobal;
		   Add083aIW	: in integer range 0 to cIWGlobal;
		   Add084aIW	: in integer range 0 to cIWGlobal;
		   Add085aIW	: in integer range 0 to cIWGlobal;
		   Add086aIW	: in integer range 0 to cIWGlobal;
		   Add087aIW	: in integer range 0 to cIWGlobal;
		   Add088aIW	: in integer range 0 to cIWGlobal;
		   Add089aIW	: in integer range 0 to cIWGlobal;
		   Add090aIW	: in integer range 0 to cIWGlobal;
		   Add091aIW	: in integer range 0 to cIWGlobal;
		   Add092aIW	: in integer range 0 to cIWGlobal;
		   Add093aIW	: in integer range 0 to cIWGlobal;
		   Add094aIW	: in integer range 0 to cIWGlobal;
		   Add095aIW	: in integer range 0 to cIWGlobal;
		   Add096aIW	: in integer range 0 to cIWGlobal;
		   Add097aIW	: in integer range 0 to cIWGlobal;
		   Add098aIW	: in integer range 0 to cIWGlobal;
		   Add099aIW	: in integer range 0 to cIWGlobal;
		   Add100aIW	: in integer range 0 to cIWGlobal;
		   Add101aIW	: in integer range 0 to cIWGlobal;
		   Add102aIW	: in integer range 0 to cIWGlobal;
		   Add103aIW	: in integer range 0 to cIWGlobal;
		   Add104aIW	: in integer range 0 to cIWGlobal;
		   Add105aIW	: in integer range 0 to cIWGlobal;
		   Add106aIW	: in integer range 0 to cIWGlobal;
		   Add107aIW	: in integer range 0 to cIWGlobal;
		   Add108aIW	: in integer range 0 to cIWGlobal;
		   Add109aIW	: in integer range 0 to cIWGlobal;
		   Add110aIW	: in integer range 0 to cIWGlobal;
		   Add111aIW	: in integer range 0 to cIWGlobal;
		   Add112aIW	: in integer range 0 to cIWGlobal;
		   Add113aIW	: in integer range 0 to cIWGlobal;
		   Add114aIW	: in integer range 0 to cIWGlobal;
		   Add115aIW	: in integer range 0 to cIWGlobal;
		   Add116aIW	: in integer range 0 to cIWGlobal;
		   Add117aIW	: in integer range 0 to cIWGlobal;
		   Add118aIW	: in integer range 0 to cIWGlobal;
		   Add119aIW	: in integer range 0 to cIWGlobal;
		   Add120aIW	: in integer range 0 to cIWGlobal;
		   Add121aIW	: in integer range 0 to cIWGlobal;
		   Add122aIW	: in integer range 0 to cIWGlobal;
		   Add123aIW	: in integer range 0 to cIWGlobal;
		   Add124aIW	: in integer range 0 to cIWGlobal;
		   Add125aIW	: in integer range 0 to cIWGlobal;
		   Add126aIW	: in integer range 0 to cIWGlobal;
		   Add127aIW	: in integer range 0 to cIWGlobal;
		   Add128aIW	: in integer range 0 to cIWGlobal;
		   Add129aIW	: in integer range 0 to cIWGlobal;
		   Add130aIW	: in integer range 0 to cIWGlobal;
		   Add131aIW	: in integer range 0 to cIWGlobal;
		   Add132aIW	: in integer range 0 to cIWGlobal;
		   Add133aIW	: in integer range 0 to cIWGlobal;
		   Add134aIW	: in integer range 0 to cIWGlobal;
		   Add135aIW	: in integer range 0 to cIWGlobal;
		   Add136aIW	: in integer range 0 to cIWGlobal;
		   Add137aIW	: in integer range 0 to cIWGlobal;
		   Add138aIW	: in integer range 0 to cIWGlobal;
		   Add139aIW	: in integer range 0 to cIWGlobal;
		   Add140aIW	: in integer range 0 to cIWGlobal;
		   Add141aIW	: in integer range 0 to cIWGlobal;
		   Add142aIW	: in integer range 0 to cIWGlobal;
		   Add143aIW	: in integer range 0 to cIWGlobal;
		   Add144aIW	: in integer range 0 to cIWGlobal;
		   Add145aIW	: in integer range 0 to cIWGlobal;
		   Add146aIW	: in integer range 0 to cIWGlobal;
		   Add147aIW	: in integer range 0 to cIWGlobal;
		   Add148aIW	: in integer range 0 to cIWGlobal;
		   Add149aIW	: in integer range 0 to cIWGlobal;
		   Add150aIW	: in integer range 0 to cIWGlobal;
		
		   Add000aFW	: in integer range 0 to cFWGlobal;
		   Add001aFW	: in integer range 0 to cFWGlobal;
		   Add002aFW	: in integer range 0 to cFWGlobal;
		   Add003aFW	: in integer range 0 to cFWGlobal;
		   Add004aFW	: in integer range 0 to cFWGlobal;
		   Add005aFW	: in integer range 0 to cFWGlobal;
		   Add006aFW	: in integer range 0 to cFWGlobal;
		   Add007aFW	: in integer range 0 to cFWGlobal;
		   Add008aFW	: in integer range 0 to cFWGlobal;
		   Add009aFW	: in integer range 0 to cFWGlobal;
		   Add010aFW	: in integer range 0 to cFWGlobal;
		   Add011aFW	: in integer range 0 to cFWGlobal;
		   Add012aFW	: in integer range 0 to cFWGlobal;
		   Add013aFW	: in integer range 0 to cFWGlobal;
		   Add014aFW	: in integer range 0 to cFWGlobal;
		   Add015aFW	: in integer range 0 to cFWGlobal;
		   Add016aFW	: in integer range 0 to cFWGlobal;
		   Add017aFW	: in integer range 0 to cFWGlobal;
		   Add018aFW	: in integer range 0 to cFWGlobal;
		   Add019aFW	: in integer range 0 to cFWGlobal;
		   Add020aFW	: in integer range 0 to cFWGlobal;
		   Add021aFW	: in integer range 0 to cFWGlobal;
		   Add022aFW	: in integer range 0 to cFWGlobal;
		   Add023aFW	: in integer range 0 to cFWGlobal;
		   Add024aFW	: in integer range 0 to cFWGlobal;
		   Add025aFW	: in integer range 0 to cFWGlobal;
		   Add026aFW	: in integer range 0 to cFWGlobal;
		   Add027aFW	: in integer range 0 to cFWGlobal;
		   Add028aFW	: in integer range 0 to cFWGlobal;
		   Add029aFW	: in integer range 0 to cFWGlobal;
		   Add030aFW	: in integer range 0 to cFWGlobal;
		   Add031aFW	: in integer range 0 to cFWGlobal;
		   Add032aFW	: in integer range 0 to cFWGlobal;
		   Add033aFW	: in integer range 0 to cFWGlobal;
		   Add034aFW	: in integer range 0 to cFWGlobal;
		   Add035aFW	: in integer range 0 to cFWGlobal;
		   Add036aFW	: in integer range 0 to cFWGlobal;
		   Add037aFW	: in integer range 0 to cFWGlobal;
		   Add038aFW	: in integer range 0 to cFWGlobal;
		   Add039aFW	: in integer range 0 to cFWGlobal;
		   Add040aFW	: in integer range 0 to cFWGlobal;
		   Add041aFW	: in integer range 0 to cFWGlobal;
		   Add042aFW	: in integer range 0 to cFWGlobal;
		   Add043aFW	: in integer range 0 to cFWGlobal;
		   Add044aFW	: in integer range 0 to cFWGlobal;
		   Add045aFW	: in integer range 0 to cFWGlobal;
		   Add046aFW	: in integer range 0 to cFWGlobal;
		   Add047aFW	: in integer range 0 to cFWGlobal;
		   Add048aFW	: in integer range 0 to cFWGlobal;
		   Add049aFW	: in integer range 0 to cFWGlobal;
		   Add050aFW	: in integer range 0 to cFWGlobal;
		   Add051aFW	: in integer range 0 to cFWGlobal;
		   Add052aFW	: in integer range 0 to cFWGlobal;
		   Add053aFW	: in integer range 0 to cFWGlobal;
		   Add054aFW	: in integer range 0 to cFWGlobal;
		   Add055aFW	: in integer range 0 to cFWGlobal;
		   Add056aFW	: in integer range 0 to cFWGlobal;
		   Add057aFW	: in integer range 0 to cFWGlobal;
		   Add058aFW	: in integer range 0 to cFWGlobal;
		   Add059aFW	: in integer range 0 to cFWGlobal;
		   Add060aFW	: in integer range 0 to cFWGlobal;
		   Add061aFW	: in integer range 0 to cFWGlobal;
		   Add062aFW	: in integer range 0 to cFWGlobal;
		   Add063aFW	: in integer range 0 to cFWGlobal;
		   Add064aFW	: in integer range 0 to cFWGlobal;
		   Add065aFW	: in integer range 0 to cFWGlobal;
		   Add066aFW	: in integer range 0 to cFWGlobal;
		   Add067aFW	: in integer range 0 to cFWGlobal;
		   Add068aFW	: in integer range 0 to cFWGlobal;
		   Add069aFW	: in integer range 0 to cFWGlobal;
		   Add070aFW	: in integer range 0 to cFWGlobal;
		   Add071aFW	: in integer range 0 to cFWGlobal;
		   Add072aFW	: in integer range 0 to cFWGlobal;
		   Add073aFW	: in integer range 0 to cFWGlobal;
		   Add074aFW	: in integer range 0 to cFWGlobal;
		   Add075aFW	: in integer range 0 to cFWGlobal;
		   Add076aFW	: in integer range 0 to cFWGlobal;
		   Add077aFW	: in integer range 0 to cFWGlobal;
		   Add078aFW	: in integer range 0 to cFWGlobal;
		   Add079aFW	: in integer range 0 to cFWGlobal;
		   Add080aFW	: in integer range 0 to cFWGlobal;
		   Add081aFW	: in integer range 0 to cFWGlobal;
		   Add082aFW	: in integer range 0 to cFWGlobal;
		   Add083aFW	: in integer range 0 to cFWGlobal;
		   Add084aFW	: in integer range 0 to cFWGlobal;
		   Add085aFW	: in integer range 0 to cFWGlobal;
		   Add086aFW	: in integer range 0 to cFWGlobal;
		   Add087aFW	: in integer range 0 to cFWGlobal;
		   Add088aFW	: in integer range 0 to cFWGlobal;
		   Add089aFW	: in integer range 0 to cFWGlobal;
		   Add090aFW	: in integer range 0 to cFWGlobal;
		   Add091aFW	: in integer range 0 to cFWGlobal;
		   Add092aFW	: in integer range 0 to cFWGlobal;
		   Add093aFW	: in integer range 0 to cFWGlobal;
		   Add094aFW	: in integer range 0 to cFWGlobal;
		   Add095aFW	: in integer range 0 to cFWGlobal;
		   Add096aFW	: in integer range 0 to cFWGlobal;
		   Add097aFW	: in integer range 0 to cFWGlobal;
		   Add098aFW	: in integer range 0 to cFWGlobal;
		   Add099aFW	: in integer range 0 to cFWGlobal;
		   Add100aFW	: in integer range 0 to cFWGlobal;
		   Add101aFW	: in integer range 0 to cFWGlobal;
		   Add102aFW	: in integer range 0 to cFWGlobal;
		   Add103aFW	: in integer range 0 to cFWGlobal;
		   Add104aFW	: in integer range 0 to cFWGlobal;
		   Add105aFW	: in integer range 0 to cFWGlobal;
		   Add106aFW	: in integer range 0 to cFWGlobal;
		   Add107aFW	: in integer range 0 to cFWGlobal;
		   Add108aFW	: in integer range 0 to cFWGlobal;
		   Add109aFW	: in integer range 0 to cFWGlobal;
		   Add110aFW	: in integer range 0 to cFWGlobal;
		   Add111aFW	: in integer range 0 to cFWGlobal;
		   Add112aFW	: in integer range 0 to cFWGlobal;
		   Add113aFW	: in integer range 0 to cFWGlobal;
		   Add114aFW	: in integer range 0 to cFWGlobal;
		   Add115aFW	: in integer range 0 to cFWGlobal;
		   Add116aFW	: in integer range 0 to cFWGlobal;
		   Add117aFW	: in integer range 0 to cFWGlobal;
		   Add118aFW	: in integer range 0 to cFWGlobal;
		   Add119aFW	: in integer range 0 to cFWGlobal;
		   Add120aFW	: in integer range 0 to cFWGlobal;
		   Add121aFW	: in integer range 0 to cFWGlobal;
		   Add122aFW	: in integer range 0 to cFWGlobal;
		   Add123aFW	: in integer range 0 to cFWGlobal;
		   Add124aFW	: in integer range 0 to cFWGlobal;
		   Add125aFW	: in integer range 0 to cFWGlobal;
		   Add126aFW	: in integer range 0 to cFWGlobal;
		   Add127aFW	: in integer range 0 to cFWGlobal;
		   Add128aFW	: in integer range 0 to cFWGlobal;
		   Add129aFW	: in integer range 0 to cFWGlobal;
		   Add130aFW	: in integer range 0 to cFWGlobal;
		   Add131aFW	: in integer range 0 to cFWGlobal;
		   Add132aFW	: in integer range 0 to cFWGlobal;
		   Add133aFW	: in integer range 0 to cFWGlobal;
		   Add134aFW	: in integer range 0 to cFWGlobal;
		   Add135aFW	: in integer range 0 to cFWGlobal;
		   Add136aFW	: in integer range 0 to cFWGlobal;
		   Add137aFW	: in integer range 0 to cFWGlobal;
		   Add138aFW	: in integer range 0 to cFWGlobal;
		   Add139aFW	: in integer range 0 to cFWGlobal;
		   Add140aFW	: in integer range 0 to cFWGlobal;
		   Add141aFW	: in integer range 0 to cFWGlobal;
		   Add142aFW	: in integer range 0 to cFWGlobal;
		   Add143aFW	: in integer range 0 to cFWGlobal;
		   Add144aFW	: in integer range 0 to cFWGlobal;
		   Add145aFW	: in integer range 0 to cFWGlobal;
		   Add146aFW	: in integer range 0 to cFWGlobal;
		   Add147aFW	: in integer range 0 to cFWGlobal;
		   Add148aFW	: in integer range 0 to cFWGlobal;
		   Add149aFW	: in integer range 0 to cFWGlobal;
		   Add150aFW	: in integer range 0 to cFWGlobal;
		   
		   Add000bIW	: in integer range 0 to cIWGlobal;
		   Add001bIW	: in integer range 0 to cIWGlobal;
		   Add002bIW	: in integer range 0 to cIWGlobal;
		   Add003bIW	: in integer range 0 to cIWGlobal;
		   Add004bIW	: in integer range 0 to cIWGlobal;
		   Add005bIW	: in integer range 0 to cIWGlobal;
		   Add006bIW	: in integer range 0 to cIWGlobal;
		   Add007bIW	: in integer range 0 to cIWGlobal;
		   Add008bIW	: in integer range 0 to cIWGlobal;
		   Add009bIW	: in integer range 0 to cIWGlobal;
		   Add010bIW	: in integer range 0 to cIWGlobal;
		   Add011bIW	: in integer range 0 to cIWGlobal;
		   Add012bIW	: in integer range 0 to cIWGlobal;
		   Add013bIW	: in integer range 0 to cIWGlobal;
		   Add014bIW	: in integer range 0 to cIWGlobal;
		   Add015bIW	: in integer range 0 to cIWGlobal;
		   Add016bIW	: in integer range 0 to cIWGlobal;
		   Add017bIW	: in integer range 0 to cIWGlobal;
		   Add018bIW	: in integer range 0 to cIWGlobal;
		   Add019bIW	: in integer range 0 to cIWGlobal;
		   Add020bIW	: in integer range 0 to cIWGlobal;
		   Add021bIW	: in integer range 0 to cIWGlobal;
		   Add022bIW	: in integer range 0 to cIWGlobal;
		   Add023bIW	: in integer range 0 to cIWGlobal;
		   Add024bIW	: in integer range 0 to cIWGlobal;
		   Add025bIW	: in integer range 0 to cIWGlobal;
		   Add026bIW	: in integer range 0 to cIWGlobal;
		   Add027bIW	: in integer range 0 to cIWGlobal;
		   Add028bIW	: in integer range 0 to cIWGlobal;
		   Add029bIW	: in integer range 0 to cIWGlobal;
		   Add030bIW	: in integer range 0 to cIWGlobal;
		   Add031bIW	: in integer range 0 to cIWGlobal;
		   Add032bIW	: in integer range 0 to cIWGlobal;
		   Add033bIW	: in integer range 0 to cIWGlobal;
		   Add034bIW	: in integer range 0 to cIWGlobal;
		   Add035bIW	: in integer range 0 to cIWGlobal;
		   Add036bIW	: in integer range 0 to cIWGlobal;
		   Add037bIW	: in integer range 0 to cIWGlobal;
		   Add038bIW	: in integer range 0 to cIWGlobal;
		   Add039bIW	: in integer range 0 to cIWGlobal;
		   Add040bIW	: in integer range 0 to cIWGlobal;
		   Add041bIW	: in integer range 0 to cIWGlobal;
		   Add042bIW	: in integer range 0 to cIWGlobal;
		   Add043bIW	: in integer range 0 to cIWGlobal;
		   Add044bIW	: in integer range 0 to cIWGlobal;
		   Add045bIW	: in integer range 0 to cIWGlobal;
		   Add046bIW	: in integer range 0 to cIWGlobal;
		   Add047bIW	: in integer range 0 to cIWGlobal;
		   Add048bIW	: in integer range 0 to cIWGlobal;
		   Add049bIW	: in integer range 0 to cIWGlobal;
		   Add050bIW	: in integer range 0 to cIWGlobal;
		   Add051bIW	: in integer range 0 to cIWGlobal;
		   Add052bIW	: in integer range 0 to cIWGlobal;
		   Add053bIW	: in integer range 0 to cIWGlobal;
		   Add054bIW	: in integer range 0 to cIWGlobal;
		   Add055bIW	: in integer range 0 to cIWGlobal;
		   Add056bIW	: in integer range 0 to cIWGlobal;
		   Add057bIW	: in integer range 0 to cIWGlobal;
		   Add058bIW	: in integer range 0 to cIWGlobal;
		   Add059bIW	: in integer range 0 to cIWGlobal;
		   Add060bIW	: in integer range 0 to cIWGlobal;
		   Add061bIW	: in integer range 0 to cIWGlobal;
		   Add062bIW	: in integer range 0 to cIWGlobal;
		   Add063bIW	: in integer range 0 to cIWGlobal;
		   Add064bIW	: in integer range 0 to cIWGlobal;
		   Add065bIW	: in integer range 0 to cIWGlobal;
		   Add066bIW	: in integer range 0 to cIWGlobal;
		   Add067bIW	: in integer range 0 to cIWGlobal;
		   Add068bIW	: in integer range 0 to cIWGlobal;
		   Add069bIW	: in integer range 0 to cIWGlobal;
		   Add070bIW	: in integer range 0 to cIWGlobal;
		   Add071bIW	: in integer range 0 to cIWGlobal;
		   Add072bIW	: in integer range 0 to cIWGlobal;
		   Add073bIW	: in integer range 0 to cIWGlobal;
		   Add074bIW	: in integer range 0 to cIWGlobal;
		   Add075bIW	: in integer range 0 to cIWGlobal;
		   Add076bIW	: in integer range 0 to cIWGlobal;
		   Add077bIW	: in integer range 0 to cIWGlobal;
		   Add078bIW	: in integer range 0 to cIWGlobal;
		   Add079bIW	: in integer range 0 to cIWGlobal;
		   Add080bIW	: in integer range 0 to cIWGlobal;
		   Add081bIW	: in integer range 0 to cIWGlobal;
		   Add082bIW	: in integer range 0 to cIWGlobal;
		   Add083bIW	: in integer range 0 to cIWGlobal;
		   Add084bIW	: in integer range 0 to cIWGlobal;
		   Add085bIW	: in integer range 0 to cIWGlobal;
		   Add086bIW	: in integer range 0 to cIWGlobal;
		   Add087bIW	: in integer range 0 to cIWGlobal;
		   Add088bIW	: in integer range 0 to cIWGlobal;
		   Add089bIW	: in integer range 0 to cIWGlobal;
		   Add090bIW	: in integer range 0 to cIWGlobal;
		   Add091bIW	: in integer range 0 to cIWGlobal;
		   Add092bIW	: in integer range 0 to cIWGlobal;
		   Add093bIW	: in integer range 0 to cIWGlobal;
		   Add094bIW	: in integer range 0 to cIWGlobal;
		   Add095bIW	: in integer range 0 to cIWGlobal;
		   Add096bIW	: in integer range 0 to cIWGlobal;
		   Add097bIW	: in integer range 0 to cIWGlobal;
		   Add098bIW	: in integer range 0 to cIWGlobal;
		   Add099bIW	: in integer range 0 to cIWGlobal;
		   Add100bIW	: in integer range 0 to cIWGlobal;
		   Add101bIW	: in integer range 0 to cIWGlobal;
		   Add102bIW	: in integer range 0 to cIWGlobal;
		   Add103bIW	: in integer range 0 to cIWGlobal;
		   Add104bIW	: in integer range 0 to cIWGlobal;
		   Add105bIW	: in integer range 0 to cIWGlobal;
		   Add106bIW	: in integer range 0 to cIWGlobal;
		   Add107bIW	: in integer range 0 to cIWGlobal;
		   Add108bIW	: in integer range 0 to cIWGlobal;
		   Add109bIW	: in integer range 0 to cIWGlobal;
		   Add110bIW	: in integer range 0 to cIWGlobal;
		   Add111bIW	: in integer range 0 to cIWGlobal;
		   Add112bIW	: in integer range 0 to cIWGlobal;
		   Add113bIW	: in integer range 0 to cIWGlobal;
		   Add114bIW	: in integer range 0 to cIWGlobal;
		   Add115bIW	: in integer range 0 to cIWGlobal;
		   Add116bIW	: in integer range 0 to cIWGlobal;
		   Add117bIW	: in integer range 0 to cIWGlobal;
		   Add118bIW	: in integer range 0 to cIWGlobal;
		   Add119bIW	: in integer range 0 to cIWGlobal;
		   Add120bIW	: in integer range 0 to cIWGlobal;
		   Add121bIW	: in integer range 0 to cIWGlobal;
		   Add122bIW	: in integer range 0 to cIWGlobal;
		   Add123bIW	: in integer range 0 to cIWGlobal;
		   Add124bIW	: in integer range 0 to cIWGlobal;
		   Add125bIW	: in integer range 0 to cIWGlobal;
		   Add126bIW	: in integer range 0 to cIWGlobal;
		   Add127bIW	: in integer range 0 to cIWGlobal;
		   Add128bIW	: in integer range 0 to cIWGlobal;
		   Add129bIW	: in integer range 0 to cIWGlobal;
		   Add130bIW	: in integer range 0 to cIWGlobal;
		   Add131bIW	: in integer range 0 to cIWGlobal;
		   Add132bIW	: in integer range 0 to cIWGlobal;
		   Add133bIW	: in integer range 0 to cIWGlobal;
		   Add134bIW	: in integer range 0 to cIWGlobal;
		   Add135bIW	: in integer range 0 to cIWGlobal;
		   Add136bIW	: in integer range 0 to cIWGlobal;
		   Add137bIW	: in integer range 0 to cIWGlobal;
		   Add138bIW	: in integer range 0 to cIWGlobal;
		   Add139bIW	: in integer range 0 to cIWGlobal;
		   Add140bIW	: in integer range 0 to cIWGlobal;
		   Add141bIW	: in integer range 0 to cIWGlobal;
		   Add142bIW	: in integer range 0 to cIWGlobal;
		   Add143bIW	: in integer range 0 to cIWGlobal;
		   Add144bIW	: in integer range 0 to cIWGlobal;
		   Add145bIW	: in integer range 0 to cIWGlobal;
		   Add146bIW	: in integer range 0 to cIWGlobal;
		   Add147bIW	: in integer range 0 to cIWGlobal;
		   Add148bIW	: in integer range 0 to cIWGlobal;
		   Add149bIW	: in integer range 0 to cIWGlobal;
		   Add150bIW	: in integer range 0 to cIWGlobal;
		 
		   Add000bFW	: in integer range 0 to cFWGlobal;
		   Add001bFW	: in integer range 0 to cFWGlobal;
		   Add002bFW	: in integer range 0 to cFWGlobal;
		   Add003bFW	: in integer range 0 to cFWGlobal;
		   Add004bFW	: in integer range 0 to cFWGlobal;
		   Add005bFW	: in integer range 0 to cFWGlobal;
		   Add006bFW	: in integer range 0 to cFWGlobal;
		   Add007bFW	: in integer range 0 to cFWGlobal;
		   Add008bFW	: in integer range 0 to cFWGlobal;
		   Add009bFW	: in integer range 0 to cFWGlobal;
		   Add010bFW	: in integer range 0 to cFWGlobal;
		   Add011bFW	: in integer range 0 to cFWGlobal;
		   Add012bFW	: in integer range 0 to cFWGlobal;
		   Add013bFW	: in integer range 0 to cFWGlobal;
		   Add014bFW	: in integer range 0 to cFWGlobal;
		   Add015bFW	: in integer range 0 to cFWGlobal;
		   Add016bFW	: in integer range 0 to cFWGlobal;
		   Add017bFW	: in integer range 0 to cFWGlobal;
		   Add018bFW	: in integer range 0 to cFWGlobal;
		   Add019bFW	: in integer range 0 to cFWGlobal;
		   Add020bFW	: in integer range 0 to cFWGlobal;
		   Add021bFW	: in integer range 0 to cFWGlobal;
		   Add022bFW	: in integer range 0 to cFWGlobal;
		   Add023bFW	: in integer range 0 to cFWGlobal;
		   Add024bFW	: in integer range 0 to cFWGlobal;
		   Add025bFW	: in integer range 0 to cFWGlobal;
		   Add026bFW	: in integer range 0 to cFWGlobal;
		   Add027bFW	: in integer range 0 to cFWGlobal;
		   Add028bFW	: in integer range 0 to cFWGlobal;
		   Add029bFW	: in integer range 0 to cFWGlobal;
		   Add030bFW	: in integer range 0 to cFWGlobal;
		   Add031bFW	: in integer range 0 to cFWGlobal;
		   Add032bFW	: in integer range 0 to cFWGlobal;
		   Add033bFW	: in integer range 0 to cFWGlobal;
		   Add034bFW	: in integer range 0 to cFWGlobal;
		   Add035bFW	: in integer range 0 to cFWGlobal;
		   Add036bFW	: in integer range 0 to cFWGlobal;
		   Add037bFW	: in integer range 0 to cFWGlobal;
		   Add038bFW	: in integer range 0 to cFWGlobal;
		   Add039bFW	: in integer range 0 to cFWGlobal;
		   Add040bFW	: in integer range 0 to cFWGlobal;
		   Add041bFW	: in integer range 0 to cFWGlobal;
		   Add042bFW	: in integer range 0 to cFWGlobal;
		   Add043bFW	: in integer range 0 to cFWGlobal;
		   Add044bFW	: in integer range 0 to cFWGlobal;
		   Add045bFW	: in integer range 0 to cFWGlobal;
		   Add046bFW	: in integer range 0 to cFWGlobal;
		   Add047bFW	: in integer range 0 to cFWGlobal;
		   Add048bFW	: in integer range 0 to cFWGlobal;
		   Add049bFW	: in integer range 0 to cFWGlobal;
		   Add050bFW	: in integer range 0 to cFWGlobal;
		   Add051bFW	: in integer range 0 to cFWGlobal;
		   Add052bFW	: in integer range 0 to cFWGlobal;
		   Add053bFW	: in integer range 0 to cFWGlobal;
		   Add054bFW	: in integer range 0 to cFWGlobal;
		   Add055bFW	: in integer range 0 to cFWGlobal;
		   Add056bFW	: in integer range 0 to cFWGlobal;
		   Add057bFW	: in integer range 0 to cFWGlobal;
		   Add058bFW	: in integer range 0 to cFWGlobal;
		   Add059bFW	: in integer range 0 to cFWGlobal;
		   Add060bFW	: in integer range 0 to cFWGlobal;
		   Add061bFW	: in integer range 0 to cFWGlobal;
		   Add062bFW	: in integer range 0 to cFWGlobal;
		   Add063bFW	: in integer range 0 to cFWGlobal;
		   Add064bFW	: in integer range 0 to cFWGlobal;
		   Add065bFW	: in integer range 0 to cFWGlobal;
		   Add066bFW	: in integer range 0 to cFWGlobal;
		   Add067bFW	: in integer range 0 to cFWGlobal;
		   Add068bFW	: in integer range 0 to cFWGlobal;
		   Add069bFW	: in integer range 0 to cFWGlobal;
		   Add070bFW	: in integer range 0 to cFWGlobal;
		   Add071bFW	: in integer range 0 to cFWGlobal;
		   Add072bFW	: in integer range 0 to cFWGlobal;
		   Add073bFW	: in integer range 0 to cFWGlobal;
		   Add074bFW	: in integer range 0 to cFWGlobal;
		   Add075bFW	: in integer range 0 to cFWGlobal;
		   Add076bFW	: in integer range 0 to cFWGlobal;
		   Add077bFW	: in integer range 0 to cFWGlobal;
		   Add078bFW	: in integer range 0 to cFWGlobal;
		   Add079bFW	: in integer range 0 to cFWGlobal;
		   Add080bFW	: in integer range 0 to cFWGlobal;
		   Add081bFW	: in integer range 0 to cFWGlobal;
		   Add082bFW	: in integer range 0 to cFWGlobal;
		   Add083bFW	: in integer range 0 to cFWGlobal;
		   Add084bFW	: in integer range 0 to cFWGlobal;
		   Add085bFW	: in integer range 0 to cFWGlobal;
		   Add086bFW	: in integer range 0 to cFWGlobal;
		   Add087bFW	: in integer range 0 to cFWGlobal;
		   Add088bFW	: in integer range 0 to cFWGlobal;
		   Add089bFW	: in integer range 0 to cFWGlobal;
		   Add090bFW	: in integer range 0 to cFWGlobal;
		   Add091bFW	: in integer range 0 to cFWGlobal;
		   Add092bFW	: in integer range 0 to cFWGlobal;
		   Add093bFW	: in integer range 0 to cFWGlobal;
		   Add094bFW	: in integer range 0 to cFWGlobal;
		   Add095bFW	: in integer range 0 to cFWGlobal;
		   Add096bFW	: in integer range 0 to cFWGlobal;
		   Add097bFW	: in integer range 0 to cFWGlobal;
		   Add098bFW	: in integer range 0 to cFWGlobal;
		   Add099bFW	: in integer range 0 to cFWGlobal;
		   Add100bFW	: in integer range 0 to cFWGlobal;
		   Add101bFW	: in integer range 0 to cFWGlobal;
		   Add102bFW	: in integer range 0 to cFWGlobal;
		   Add103bFW	: in integer range 0 to cFWGlobal;
		   Add104bFW	: in integer range 0 to cFWGlobal;
		   Add105bFW	: in integer range 0 to cFWGlobal;
		   Add106bFW	: in integer range 0 to cFWGlobal;
		   Add107bFW	: in integer range 0 to cFWGlobal;
		   Add108bFW	: in integer range 0 to cFWGlobal;
		   Add109bFW	: in integer range 0 to cFWGlobal;
		   Add110bFW	: in integer range 0 to cFWGlobal;
		   Add111bFW	: in integer range 0 to cFWGlobal;
		   Add112bFW	: in integer range 0 to cFWGlobal;
		   Add113bFW	: in integer range 0 to cFWGlobal;
		   Add114bFW	: in integer range 0 to cFWGlobal;
		   Add115bFW	: in integer range 0 to cFWGlobal;
		   Add116bFW	: in integer range 0 to cFWGlobal;
		   Add117bFW	: in integer range 0 to cFWGlobal;
		   Add118bFW	: in integer range 0 to cFWGlobal;
		   Add119bFW	: in integer range 0 to cFWGlobal;
		   Add120bFW	: in integer range 0 to cFWGlobal;
		   Add121bFW	: in integer range 0 to cFWGlobal;
		   Add122bFW	: in integer range 0 to cFWGlobal;
		   Add123bFW	: in integer range 0 to cFWGlobal;
		   Add124bFW	: in integer range 0 to cFWGlobal;
		   Add125bFW	: in integer range 0 to cFWGlobal;
		   Add126bFW	: in integer range 0 to cFWGlobal;
		   Add127bFW	: in integer range 0 to cFWGlobal;
		   Add128bFW	: in integer range 0 to cFWGlobal;
		   Add129bFW	: in integer range 0 to cFWGlobal;
		   Add130bFW	: in integer range 0 to cFWGlobal;
		   Add131bFW	: in integer range 0 to cFWGlobal;
		   Add132bFW	: in integer range 0 to cFWGlobal;
		   Add133bFW	: in integer range 0 to cFWGlobal;
		   Add134bFW	: in integer range 0 to cFWGlobal;
		   Add135bFW	: in integer range 0 to cFWGlobal;
		   Add136bFW	: in integer range 0 to cFWGlobal;
		   Add137bFW	: in integer range 0 to cFWGlobal;
		   Add138bFW	: in integer range 0 to cFWGlobal;
		   Add139bFW	: in integer range 0 to cFWGlobal;
		   Add140bFW	: in integer range 0 to cFWGlobal;
		   Add141bFW	: in integer range 0 to cFWGlobal;
		   Add142bFW	: in integer range 0 to cFWGlobal;
		   Add143bFW	: in integer range 0 to cFWGlobal;
		   Add144bFW	: in integer range 0 to cFWGlobal;
		   Add145bFW	: in integer range 0 to cFWGlobal;
		   Add146bFW	: in integer range 0 to cFWGlobal;
		   Add147bFW	: in integer range 0 to cFWGlobal;
		   Add148bFW	: in integer range 0 to cFWGlobal;
		   Add149bFW	: in integer range 0 to cFWGlobal;
		   Add150bFW	: in integer range 0 to cFWGlobal;
		   
		   
		   
		   Mult000aIW	: in integer range 0 to cIWGlobal;
		   Mult001aIW	: in integer range 0 to cIWGlobal;
		   Mult002aIW	: in integer range 0 to cIWGlobal;
		   Mult003aIW	: in integer range 0 to cIWGlobal;
		   Mult004aIW	: in integer range 0 to cIWGlobal;
		   Mult005aIW	: in integer range 0 to cIWGlobal;
		   Mult006aIW	: in integer range 0 to cIWGlobal;
		   Mult007aIW	: in integer range 0 to cIWGlobal;
		   Mult008aIW	: in integer range 0 to cIWGlobal;
		   Mult009aIW	: in integer range 0 to cIWGlobal;
		   Mult010aIW	: in integer range 0 to cIWGlobal;
		   Mult011aIW	: in integer range 0 to cIWGlobal;
		   Mult012aIW	: in integer range 0 to cIWGlobal;
		   Mult013aIW	: in integer range 0 to cIWGlobal;
		   Mult014aIW	: in integer range 0 to cIWGlobal;
		   Mult015aIW	: in integer range 0 to cIWGlobal;
		   Mult016aIW	: in integer range 0 to cIWGlobal;
		   Mult017aIW	: in integer range 0 to cIWGlobal;
		   Mult018aIW	: in integer range 0 to cIWGlobal;
		   Mult019aIW	: in integer range 0 to cIWGlobal;
		   Mult020aIW	: in integer range 0 to cIWGlobal;
		   Mult021aIW	: in integer range 0 to cIWGlobal;
		   Mult022aIW	: in integer range 0 to cIWGlobal;
		   Mult023aIW	: in integer range 0 to cIWGlobal;
		   Mult024aIW	: in integer range 0 to cIWGlobal;
		   Mult025aIW	: in integer range 0 to cIWGlobal;
		   Mult026aIW	: in integer range 0 to cIWGlobal;
		   Mult027aIW	: in integer range 0 to cIWGlobal;
		   Mult028aIW	: in integer range 0 to cIWGlobal;
		   Mult029aIW	: in integer range 0 to cIWGlobal;
		   Mult030aIW	: in integer range 0 to cIWGlobal;
		   Mult031aIW	: in integer range 0 to cIWGlobal;
		   Mult032aIW	: in integer range 0 to cIWGlobal;
		   Mult033aIW	: in integer range 0 to cIWGlobal;
		   Mult034aIW	: in integer range 0 to cIWGlobal;
		   Mult035aIW	: in integer range 0 to cIWGlobal;
		   Mult036aIW	: in integer range 0 to cIWGlobal;
		   Mult037aIW	: in integer range 0 to cIWGlobal;
		   Mult038aIW	: in integer range 0 to cIWGlobal;
		   Mult039aIW	: in integer range 0 to cIWGlobal;
		   Mult040aIW	: in integer range 0 to cIWGlobal;
		   Mult041aIW	: in integer range 0 to cIWGlobal;
		   Mult042aIW	: in integer range 0 to cIWGlobal;
		   Mult043aIW	: in integer range 0 to cIWGlobal;
		   Mult044aIW	: in integer range 0 to cIWGlobal;
		   Mult045aIW	: in integer range 0 to cIWGlobal;
		   Mult046aIW	: in integer range 0 to cIWGlobal;
		   Mult047aIW	: in integer range 0 to cIWGlobal;
		   Mult048aIW	: in integer range 0 to cIWGlobal;
		   Mult049aIW	: in integer range 0 to cIWGlobal;
		   Mult050aIW	: in integer range 0 to cIWGlobal;
		   Mult051aIW	: in integer range 0 to cIWGlobal;
		   Mult052aIW	: in integer range 0 to cIWGlobal;
		   Mult053aIW	: in integer range 0 to cIWGlobal;
		   Mult054aIW	: in integer range 0 to cIWGlobal;
		   Mult055aIW	: in integer range 0 to cIWGlobal;
		   Mult056aIW	: in integer range 0 to cIWGlobal;
		   Mult057aIW	: in integer range 0 to cIWGlobal;
		   Mult058aIW	: in integer range 0 to cIWGlobal;
		   Mult059aIW	: in integer range 0 to cIWGlobal;
		   Mult060aIW	: in integer range 0 to cIWGlobal;
		   Mult061aIW	: in integer range 0 to cIWGlobal;
		   Mult062aIW	: in integer range 0 to cIWGlobal;
		   Mult063aIW	: in integer range 0 to cIWGlobal;
		   Mult064aIW	: in integer range 0 to cIWGlobal;
		   Mult065aIW	: in integer range 0 to cIWGlobal;
		   Mult066aIW	: in integer range 0 to cIWGlobal;
		   Mult067aIW	: in integer range 0 to cIWGlobal;
		   Mult068aIW	: in integer range 0 to cIWGlobal;
		   Mult069aIW	: in integer range 0 to cIWGlobal;
		   Mult070aIW	: in integer range 0 to cIWGlobal;
		   Mult071aIW	: in integer range 0 to cIWGlobal;
		   Mult072aIW	: in integer range 0 to cIWGlobal;
		   Mult073aIW	: in integer range 0 to cIWGlobal;
		   Mult074aIW	: in integer range 0 to cIWGlobal;
		   Mult075aIW	: in integer range 0 to cIWGlobal;
		   Mult076aIW	: in integer range 0 to cIWGlobal;
		   Mult077aIW	: in integer range 0 to cIWGlobal;
		   Mult078aIW	: in integer range 0 to cIWGlobal;
		   Mult079aIW	: in integer range 0 to cIWGlobal;
		   Mult080aIW	: in integer range 0 to cIWGlobal;
		   Mult081aIW	: in integer range 0 to cIWGlobal;
		   Mult082aIW	: in integer range 0 to cIWGlobal;
		   Mult083aIW	: in integer range 0 to cIWGlobal;
		   Mult084aIW	: in integer range 0 to cIWGlobal;
		   Mult085aIW	: in integer range 0 to cIWGlobal;
		   Mult086aIW	: in integer range 0 to cIWGlobal;
		   Mult087aIW	: in integer range 0 to cIWGlobal;
		   Mult088aIW	: in integer range 0 to cIWGlobal;
		   Mult089aIW	: in integer range 0 to cIWGlobal;
		   Mult090aIW	: in integer range 0 to cIWGlobal;
		   Mult091aIW	: in integer range 0 to cIWGlobal;
		   Mult092aIW	: in integer range 0 to cIWGlobal;
		   Mult093aIW	: in integer range 0 to cIWGlobal;
		   Mult094aIW	: in integer range 0 to cIWGlobal;
		   Mult095aIW	: in integer range 0 to cIWGlobal;
		   Mult096aIW	: in integer range 0 to cIWGlobal;
		   Mult097aIW	: in integer range 0 to cIWGlobal;
		   Mult098aIW	: in integer range 0 to cIWGlobal;
		   Mult099aIW	: in integer range 0 to cIWGlobal;
		   Mult100aIW	: in integer range 0 to cIWGlobal;
		   Mult101aIW	: in integer range 0 to cIWGlobal;
		   Mult102aIW	: in integer range 0 to cIWGlobal;
		   Mult103aIW	: in integer range 0 to cIWGlobal;
		   Mult104aIW	: in integer range 0 to cIWGlobal;
		   Mult105aIW	: in integer range 0 to cIWGlobal;
		   Mult106aIW	: in integer range 0 to cIWGlobal;
		   Mult107aIW	: in integer range 0 to cIWGlobal;
		   Mult108aIW	: in integer range 0 to cIWGlobal;
		   Mult109aIW	: in integer range 0 to cIWGlobal;
		   Mult110aIW	: in integer range 0 to cIWGlobal;
		   Mult111aIW	: in integer range 0 to cIWGlobal;
		   Mult112aIW	: in integer range 0 to cIWGlobal;
		   Mult113aIW	: in integer range 0 to cIWGlobal;
		   Mult114aIW	: in integer range 0 to cIWGlobal;
		   Mult115aIW	: in integer range 0 to cIWGlobal;
		   Mult116aIW	: in integer range 0 to cIWGlobal;
		   Mult117aIW	: in integer range 0 to cIWGlobal;
		   Mult118aIW	: in integer range 0 to cIWGlobal;
		   Mult119aIW	: in integer range 0 to cIWGlobal;
		   Mult120aIW	: in integer range 0 to cIWGlobal;
		   Mult121aIW	: in integer range 0 to cIWGlobal;
		   Mult122aIW	: in integer range 0 to cIWGlobal;
		   Mult123aIW	: in integer range 0 to cIWGlobal;
		   Mult124aIW	: in integer range 0 to cIWGlobal;
		   Mult125aIW	: in integer range 0 to cIWGlobal;
		   Mult126aIW	: in integer range 0 to cIWGlobal;
		   Mult127aIW	: in integer range 0 to cIWGlobal;
		   Mult128aIW	: in integer range 0 to cIWGlobal;
		   Mult129aIW	: in integer range 0 to cIWGlobal;
		   Mult130aIW	: in integer range 0 to cIWGlobal;
		   Mult131aIW	: in integer range 0 to cIWGlobal;
		   Mult132aIW	: in integer range 0 to cIWGlobal;
		   Mult133aIW	: in integer range 0 to cIWGlobal;
		   Mult134aIW	: in integer range 0 to cIWGlobal;
		   Mult135aIW	: in integer range 0 to cIWGlobal;
		   Mult136aIW	: in integer range 0 to cIWGlobal;
		   Mult137aIW	: in integer range 0 to cIWGlobal;
		   Mult138aIW	: in integer range 0 to cIWGlobal;
		   Mult139aIW	: in integer range 0 to cIWGlobal;
		   Mult140aIW	: in integer range 0 to cIWGlobal;
		   Mult141aIW	: in integer range 0 to cIWGlobal;
		   Mult142aIW	: in integer range 0 to cIWGlobal;
		   Mult143aIW	: in integer range 0 to cIWGlobal;
		   Mult144aIW	: in integer range 0 to cIWGlobal;
		   Mult145aIW	: in integer range 0 to cIWGlobal;
		   Mult146aIW	: in integer range 0 to cIWGlobal;
		   Mult147aIW	: in integer range 0 to cIWGlobal;
		   Mult148aIW	: in integer range 0 to cIWGlobal;
		   Mult149aIW	: in integer range 0 to cIWGlobal;
		   Mult150aIW	: in integer range 0 to cIWGlobal;
		
		   Mult000aFW	: in integer range 0 to cFWGlobal;
		   Mult001aFW	: in integer range 0 to cFWGlobal;
		   Mult002aFW	: in integer range 0 to cFWGlobal;
		   Mult003aFW	: in integer range 0 to cFWGlobal;
		   Mult004aFW	: in integer range 0 to cFWGlobal;
		   Mult005aFW	: in integer range 0 to cFWGlobal;
		   Mult006aFW	: in integer range 0 to cFWGlobal;
		   Mult007aFW	: in integer range 0 to cFWGlobal;
		   Mult008aFW	: in integer range 0 to cFWGlobal;
		   Mult009aFW	: in integer range 0 to cFWGlobal;
		   Mult010aFW	: in integer range 0 to cFWGlobal;
		   Mult011aFW	: in integer range 0 to cFWGlobal;
		   Mult012aFW	: in integer range 0 to cFWGlobal;
		   Mult013aFW	: in integer range 0 to cFWGlobal;
		   Mult014aFW	: in integer range 0 to cFWGlobal;
		   Mult015aFW	: in integer range 0 to cFWGlobal;
		   Mult016aFW	: in integer range 0 to cFWGlobal;
		   Mult017aFW	: in integer range 0 to cFWGlobal;
		   Mult018aFW	: in integer range 0 to cFWGlobal;
		   Mult019aFW	: in integer range 0 to cFWGlobal;
		   Mult020aFW	: in integer range 0 to cFWGlobal;
		   Mult021aFW	: in integer range 0 to cFWGlobal;
		   Mult022aFW	: in integer range 0 to cFWGlobal;
		   Mult023aFW	: in integer range 0 to cFWGlobal;
		   Mult024aFW	: in integer range 0 to cFWGlobal;
		   Mult025aFW	: in integer range 0 to cFWGlobal;
		   Mult026aFW	: in integer range 0 to cFWGlobal;
		   Mult027aFW	: in integer range 0 to cFWGlobal;
		   Mult028aFW	: in integer range 0 to cFWGlobal;
		   Mult029aFW	: in integer range 0 to cFWGlobal;
		   Mult030aFW	: in integer range 0 to cFWGlobal;
		   Mult031aFW	: in integer range 0 to cFWGlobal;
		   Mult032aFW	: in integer range 0 to cFWGlobal;
		   Mult033aFW	: in integer range 0 to cFWGlobal;
		   Mult034aFW	: in integer range 0 to cFWGlobal;
		   Mult035aFW	: in integer range 0 to cFWGlobal;
		   Mult036aFW	: in integer range 0 to cFWGlobal;
		   Mult037aFW	: in integer range 0 to cFWGlobal;
		   Mult038aFW	: in integer range 0 to cFWGlobal;
		   Mult039aFW	: in integer range 0 to cFWGlobal;
		   Mult040aFW	: in integer range 0 to cFWGlobal;
		   Mult041aFW	: in integer range 0 to cFWGlobal;
		   Mult042aFW	: in integer range 0 to cFWGlobal;
		   Mult043aFW	: in integer range 0 to cFWGlobal;
		   Mult044aFW	: in integer range 0 to cFWGlobal;
		   Mult045aFW	: in integer range 0 to cFWGlobal;
		   Mult046aFW	: in integer range 0 to cFWGlobal;
		   Mult047aFW	: in integer range 0 to cFWGlobal;
		   Mult048aFW	: in integer range 0 to cFWGlobal;
		   Mult049aFW	: in integer range 0 to cFWGlobal;
		   Mult050aFW	: in integer range 0 to cFWGlobal;
		   Mult051aFW	: in integer range 0 to cFWGlobal;
		   Mult052aFW	: in integer range 0 to cFWGlobal;
		   Mult053aFW	: in integer range 0 to cFWGlobal;
		   Mult054aFW	: in integer range 0 to cFWGlobal;
		   Mult055aFW	: in integer range 0 to cFWGlobal;
		   Mult056aFW	: in integer range 0 to cFWGlobal;
		   Mult057aFW	: in integer range 0 to cFWGlobal;
		   Mult058aFW	: in integer range 0 to cFWGlobal;
		   Mult059aFW	: in integer range 0 to cFWGlobal;
		   Mult060aFW	: in integer range 0 to cFWGlobal;
		   Mult061aFW	: in integer range 0 to cFWGlobal;
		   Mult062aFW	: in integer range 0 to cFWGlobal;
		   Mult063aFW	: in integer range 0 to cFWGlobal;
		   Mult064aFW	: in integer range 0 to cFWGlobal;
		   Mult065aFW	: in integer range 0 to cFWGlobal;
		   Mult066aFW	: in integer range 0 to cFWGlobal;
		   Mult067aFW	: in integer range 0 to cFWGlobal;
		   Mult068aFW	: in integer range 0 to cFWGlobal;
		   Mult069aFW	: in integer range 0 to cFWGlobal;
		   Mult070aFW	: in integer range 0 to cFWGlobal;
		   Mult071aFW	: in integer range 0 to cFWGlobal;
		   Mult072aFW	: in integer range 0 to cFWGlobal;
		   Mult073aFW	: in integer range 0 to cFWGlobal;
		   Mult074aFW	: in integer range 0 to cFWGlobal;
		   Mult075aFW	: in integer range 0 to cFWGlobal;
		   Mult076aFW	: in integer range 0 to cFWGlobal;
		   Mult077aFW	: in integer range 0 to cFWGlobal;
		   Mult078aFW	: in integer range 0 to cFWGlobal;
		   Mult079aFW	: in integer range 0 to cFWGlobal;
		   Mult080aFW	: in integer range 0 to cFWGlobal;
		   Mult081aFW	: in integer range 0 to cFWGlobal;
		   Mult082aFW	: in integer range 0 to cFWGlobal;
		   Mult083aFW	: in integer range 0 to cFWGlobal;
		   Mult084aFW	: in integer range 0 to cFWGlobal;
		   Mult085aFW	: in integer range 0 to cFWGlobal;
		   Mult086aFW	: in integer range 0 to cFWGlobal;
		   Mult087aFW	: in integer range 0 to cFWGlobal;
		   Mult088aFW	: in integer range 0 to cFWGlobal;
		   Mult089aFW	: in integer range 0 to cFWGlobal;
		   Mult090aFW	: in integer range 0 to cFWGlobal;
		   Mult091aFW	: in integer range 0 to cFWGlobal;
		   Mult092aFW	: in integer range 0 to cFWGlobal;
		   Mult093aFW	: in integer range 0 to cFWGlobal;
		   Mult094aFW	: in integer range 0 to cFWGlobal;
		   Mult095aFW	: in integer range 0 to cFWGlobal;
		   Mult096aFW	: in integer range 0 to cFWGlobal;
		   Mult097aFW	: in integer range 0 to cFWGlobal;
		   Mult098aFW	: in integer range 0 to cFWGlobal;
		   Mult099aFW	: in integer range 0 to cFWGlobal;
		   Mult100aFW	: in integer range 0 to cFWGlobal;
		   Mult101aFW	: in integer range 0 to cFWGlobal;
		   Mult102aFW	: in integer range 0 to cFWGlobal;
		   Mult103aFW	: in integer range 0 to cFWGlobal;
		   Mult104aFW	: in integer range 0 to cFWGlobal;
		   Mult105aFW	: in integer range 0 to cFWGlobal;
		   Mult106aFW	: in integer range 0 to cFWGlobal;
		   Mult107aFW	: in integer range 0 to cFWGlobal;
		   Mult108aFW	: in integer range 0 to cFWGlobal;
		   Mult109aFW	: in integer range 0 to cFWGlobal;
		   Mult110aFW	: in integer range 0 to cFWGlobal;
		   Mult111aFW	: in integer range 0 to cFWGlobal;
		   Mult112aFW	: in integer range 0 to cFWGlobal;
		   Mult113aFW	: in integer range 0 to cFWGlobal;
		   Mult114aFW	: in integer range 0 to cFWGlobal;
		   Mult115aFW	: in integer range 0 to cFWGlobal;
		   Mult116aFW	: in integer range 0 to cFWGlobal;
		   Mult117aFW	: in integer range 0 to cFWGlobal;
		   Mult118aFW	: in integer range 0 to cFWGlobal;
		   Mult119aFW	: in integer range 0 to cFWGlobal;
		   Mult120aFW	: in integer range 0 to cFWGlobal;
		   Mult121aFW	: in integer range 0 to cFWGlobal;
		   Mult122aFW	: in integer range 0 to cFWGlobal;
		   Mult123aFW	: in integer range 0 to cFWGlobal;
		   Mult124aFW	: in integer range 0 to cFWGlobal;
		   Mult125aFW	: in integer range 0 to cFWGlobal;
		   Mult126aFW	: in integer range 0 to cFWGlobal;
		   Mult127aFW	: in integer range 0 to cFWGlobal;
		   Mult128aFW	: in integer range 0 to cFWGlobal;
		   Mult129aFW	: in integer range 0 to cFWGlobal;
		   Mult130aFW	: in integer range 0 to cFWGlobal;
		   Mult131aFW	: in integer range 0 to cFWGlobal;
		   Mult132aFW	: in integer range 0 to cFWGlobal;
		   Mult133aFW	: in integer range 0 to cFWGlobal;
		   Mult134aFW	: in integer range 0 to cFWGlobal;
		   Mult135aFW	: in integer range 0 to cFWGlobal;
		   Mult136aFW	: in integer range 0 to cFWGlobal;
		   Mult137aFW	: in integer range 0 to cFWGlobal;
		   Mult138aFW	: in integer range 0 to cFWGlobal;
		   Mult139aFW	: in integer range 0 to cFWGlobal;
		   Mult140aFW	: in integer range 0 to cFWGlobal;
		   Mult141aFW	: in integer range 0 to cFWGlobal;
		   Mult142aFW	: in integer range 0 to cFWGlobal;
		   Mult143aFW	: in integer range 0 to cFWGlobal;
		   Mult144aFW	: in integer range 0 to cFWGlobal;
		   Mult145aFW	: in integer range 0 to cFWGlobal;
		   Mult146aFW	: in integer range 0 to cFWGlobal;
		   Mult147aFW	: in integer range 0 to cFWGlobal;
		   Mult148aFW	: in integer range 0 to cFWGlobal;
		   Mult149aFW	: in integer range 0 to cFWGlobal;
		   Mult150aFW	: in integer range 0 to cFWGlobal;
		   
		   Mult000bIW	: in integer range 0 to cIWGlobal;
		   Mult001bIW	: in integer range 0 to cIWGlobal;
		   Mult002bIW	: in integer range 0 to cIWGlobal;
		   Mult003bIW	: in integer range 0 to cIWGlobal;
		   Mult004bIW	: in integer range 0 to cIWGlobal;
		   Mult005bIW	: in integer range 0 to cIWGlobal;
		   Mult006bIW	: in integer range 0 to cIWGlobal;
		   Mult007bIW	: in integer range 0 to cIWGlobal;
		   Mult008bIW	: in integer range 0 to cIWGlobal;
		   Mult009bIW	: in integer range 0 to cIWGlobal;
		   Mult010bIW	: in integer range 0 to cIWGlobal;
		   Mult011bIW	: in integer range 0 to cIWGlobal;
		   Mult012bIW	: in integer range 0 to cIWGlobal;
		   Mult013bIW	: in integer range 0 to cIWGlobal;
		   Mult014bIW	: in integer range 0 to cIWGlobal;
		   Mult015bIW	: in integer range 0 to cIWGlobal;
		   Mult016bIW	: in integer range 0 to cIWGlobal;
		   Mult017bIW	: in integer range 0 to cIWGlobal;
		   Mult018bIW	: in integer range 0 to cIWGlobal;
		   Mult019bIW	: in integer range 0 to cIWGlobal;
		   Mult020bIW	: in integer range 0 to cIWGlobal;
		   Mult021bIW	: in integer range 0 to cIWGlobal;
		   Mult022bIW	: in integer range 0 to cIWGlobal;
		   Mult023bIW	: in integer range 0 to cIWGlobal;
		   Mult024bIW	: in integer range 0 to cIWGlobal;
		   Mult025bIW	: in integer range 0 to cIWGlobal;
		   Mult026bIW	: in integer range 0 to cIWGlobal;
		   Mult027bIW	: in integer range 0 to cIWGlobal;
		   Mult028bIW	: in integer range 0 to cIWGlobal;
		   Mult029bIW	: in integer range 0 to cIWGlobal;
		   Mult030bIW	: in integer range 0 to cIWGlobal;
		   Mult031bIW	: in integer range 0 to cIWGlobal;
		   Mult032bIW	: in integer range 0 to cIWGlobal;
		   Mult033bIW	: in integer range 0 to cIWGlobal;
		   Mult034bIW	: in integer range 0 to cIWGlobal;
		   Mult035bIW	: in integer range 0 to cIWGlobal;
		   Mult036bIW	: in integer range 0 to cIWGlobal;
		   Mult037bIW	: in integer range 0 to cIWGlobal;
		   Mult038bIW	: in integer range 0 to cIWGlobal;
		   Mult039bIW	: in integer range 0 to cIWGlobal;
		   Mult040bIW	: in integer range 0 to cIWGlobal;
		   Mult041bIW	: in integer range 0 to cIWGlobal;
		   Mult042bIW	: in integer range 0 to cIWGlobal;
		   Mult043bIW	: in integer range 0 to cIWGlobal;
		   Mult044bIW	: in integer range 0 to cIWGlobal;
		   Mult045bIW	: in integer range 0 to cIWGlobal;
		   Mult046bIW	: in integer range 0 to cIWGlobal;
		   Mult047bIW	: in integer range 0 to cIWGlobal;
		   Mult048bIW	: in integer range 0 to cIWGlobal;
		   Mult049bIW	: in integer range 0 to cIWGlobal;
		   Mult050bIW	: in integer range 0 to cIWGlobal;
		   Mult051bIW	: in integer range 0 to cIWGlobal;
		   Mult052bIW	: in integer range 0 to cIWGlobal;
		   Mult053bIW	: in integer range 0 to cIWGlobal;
		   Mult054bIW	: in integer range 0 to cIWGlobal;
		   Mult055bIW	: in integer range 0 to cIWGlobal;
		   Mult056bIW	: in integer range 0 to cIWGlobal;
		   Mult057bIW	: in integer range 0 to cIWGlobal;
		   Mult058bIW	: in integer range 0 to cIWGlobal;
		   Mult059bIW	: in integer range 0 to cIWGlobal;
		   Mult060bIW	: in integer range 0 to cIWGlobal;
		   Mult061bIW	: in integer range 0 to cIWGlobal;
		   Mult062bIW	: in integer range 0 to cIWGlobal;
		   Mult063bIW	: in integer range 0 to cIWGlobal;
		   Mult064bIW	: in integer range 0 to cIWGlobal;
		   Mult065bIW	: in integer range 0 to cIWGlobal;
		   Mult066bIW	: in integer range 0 to cIWGlobal;
		   Mult067bIW	: in integer range 0 to cIWGlobal;
		   Mult068bIW	: in integer range 0 to cIWGlobal;
		   Mult069bIW	: in integer range 0 to cIWGlobal;
		   Mult070bIW	: in integer range 0 to cIWGlobal;
		   Mult071bIW	: in integer range 0 to cIWGlobal;
		   Mult072bIW	: in integer range 0 to cIWGlobal;
		   Mult073bIW	: in integer range 0 to cIWGlobal;
		   Mult074bIW	: in integer range 0 to cIWGlobal;
		   Mult075bIW	: in integer range 0 to cIWGlobal;
		   Mult076bIW	: in integer range 0 to cIWGlobal;
		   Mult077bIW	: in integer range 0 to cIWGlobal;
		   Mult078bIW	: in integer range 0 to cIWGlobal;
		   Mult079bIW	: in integer range 0 to cIWGlobal;
		   Mult080bIW	: in integer range 0 to cIWGlobal;
		   Mult081bIW	: in integer range 0 to cIWGlobal;
		   Mult082bIW	: in integer range 0 to cIWGlobal;
		   Mult083bIW	: in integer range 0 to cIWGlobal;
		   Mult084bIW	: in integer range 0 to cIWGlobal;
		   Mult085bIW	: in integer range 0 to cIWGlobal;
		   Mult086bIW	: in integer range 0 to cIWGlobal;
		   Mult087bIW	: in integer range 0 to cIWGlobal;
		   Mult088bIW	: in integer range 0 to cIWGlobal;
		   Mult089bIW	: in integer range 0 to cIWGlobal;
		   Mult090bIW	: in integer range 0 to cIWGlobal;
		   Mult091bIW	: in integer range 0 to cIWGlobal;
		   Mult092bIW	: in integer range 0 to cIWGlobal;
		   Mult093bIW	: in integer range 0 to cIWGlobal;
		   Mult094bIW	: in integer range 0 to cIWGlobal;
		   Mult095bIW	: in integer range 0 to cIWGlobal;
		   Mult096bIW	: in integer range 0 to cIWGlobal;
		   Mult097bIW	: in integer range 0 to cIWGlobal;
		   Mult098bIW	: in integer range 0 to cIWGlobal;
		   Mult099bIW	: in integer range 0 to cIWGlobal;
		   Mult100bIW	: in integer range 0 to cIWGlobal;
		   Mult101bIW	: in integer range 0 to cIWGlobal;
		   Mult102bIW	: in integer range 0 to cIWGlobal;
		   Mult103bIW	: in integer range 0 to cIWGlobal;
		   Mult104bIW	: in integer range 0 to cIWGlobal;
		   Mult105bIW	: in integer range 0 to cIWGlobal;
		   Mult106bIW	: in integer range 0 to cIWGlobal;
		   Mult107bIW	: in integer range 0 to cIWGlobal;
		   Mult108bIW	: in integer range 0 to cIWGlobal;
		   Mult109bIW	: in integer range 0 to cIWGlobal;
		   Mult110bIW	: in integer range 0 to cIWGlobal;
		   Mult111bIW	: in integer range 0 to cIWGlobal;
		   Mult112bIW	: in integer range 0 to cIWGlobal;
		   Mult113bIW	: in integer range 0 to cIWGlobal;
		   Mult114bIW	: in integer range 0 to cIWGlobal;
		   Mult115bIW	: in integer range 0 to cIWGlobal;
		   Mult116bIW	: in integer range 0 to cIWGlobal;
		   Mult117bIW	: in integer range 0 to cIWGlobal;
		   Mult118bIW	: in integer range 0 to cIWGlobal;
		   Mult119bIW	: in integer range 0 to cIWGlobal;
		   Mult120bIW	: in integer range 0 to cIWGlobal;
		   Mult121bIW	: in integer range 0 to cIWGlobal;
		   Mult122bIW	: in integer range 0 to cIWGlobal;
		   Mult123bIW	: in integer range 0 to cIWGlobal;
		   Mult124bIW	: in integer range 0 to cIWGlobal;
		   Mult125bIW	: in integer range 0 to cIWGlobal;
		   Mult126bIW	: in integer range 0 to cIWGlobal;
		   Mult127bIW	: in integer range 0 to cIWGlobal;
		   Mult128bIW	: in integer range 0 to cIWGlobal;
		   Mult129bIW	: in integer range 0 to cIWGlobal;
		   Mult130bIW	: in integer range 0 to cIWGlobal;
		   Mult131bIW	: in integer range 0 to cIWGlobal;
		   Mult132bIW	: in integer range 0 to cIWGlobal;
		   Mult133bIW	: in integer range 0 to cIWGlobal;
		   Mult134bIW	: in integer range 0 to cIWGlobal;
		   Mult135bIW	: in integer range 0 to cIWGlobal;
		   Mult136bIW	: in integer range 0 to cIWGlobal;
		   Mult137bIW	: in integer range 0 to cIWGlobal;
		   Mult138bIW	: in integer range 0 to cIWGlobal;
		   Mult139bIW	: in integer range 0 to cIWGlobal;
		   Mult140bIW	: in integer range 0 to cIWGlobal;
		   Mult141bIW	: in integer range 0 to cIWGlobal;
		   Mult142bIW	: in integer range 0 to cIWGlobal;
		   Mult143bIW	: in integer range 0 to cIWGlobal;
		   Mult144bIW	: in integer range 0 to cIWGlobal;
		   Mult145bIW	: in integer range 0 to cIWGlobal;
		   Mult146bIW	: in integer range 0 to cIWGlobal;
		   Mult147bIW	: in integer range 0 to cIWGlobal;
		   Mult148bIW	: in integer range 0 to cIWGlobal;
		   Mult149bIW	: in integer range 0 to cIWGlobal;
		   Mult150bIW	: in integer range 0 to cIWGlobal;
		 
		   Mult000bFW	: in integer range 0 to cFWGlobal;
		   Mult001bFW	: in integer range 0 to cFWGlobal;
		   Mult002bFW	: in integer range 0 to cFWGlobal;
		   Mult003bFW	: in integer range 0 to cFWGlobal;
		   Mult004bFW	: in integer range 0 to cFWGlobal;
		   Mult005bFW	: in integer range 0 to cFWGlobal;
		   Mult006bFW	: in integer range 0 to cFWGlobal;
		   Mult007bFW	: in integer range 0 to cFWGlobal;
		   Mult008bFW	: in integer range 0 to cFWGlobal;
		   Mult009bFW	: in integer range 0 to cFWGlobal;
		   Mult010bFW	: in integer range 0 to cFWGlobal;
		   Mult011bFW	: in integer range 0 to cFWGlobal;
		   Mult012bFW	: in integer range 0 to cFWGlobal;
		   Mult013bFW	: in integer range 0 to cFWGlobal;
		   Mult014bFW	: in integer range 0 to cFWGlobal;
		   Mult015bFW	: in integer range 0 to cFWGlobal;
		   Mult016bFW	: in integer range 0 to cFWGlobal;
		   Mult017bFW	: in integer range 0 to cFWGlobal;
		   Mult018bFW	: in integer range 0 to cFWGlobal;
		   Mult019bFW	: in integer range 0 to cFWGlobal;
		   Mult020bFW	: in integer range 0 to cFWGlobal;
		   Mult021bFW	: in integer range 0 to cFWGlobal;
		   Mult022bFW	: in integer range 0 to cFWGlobal;
		   Mult023bFW	: in integer range 0 to cFWGlobal;
		   Mult024bFW	: in integer range 0 to cFWGlobal;
		   Mult025bFW	: in integer range 0 to cFWGlobal;
		   Mult026bFW	: in integer range 0 to cFWGlobal;
		   Mult027bFW	: in integer range 0 to cFWGlobal;
		   Mult028bFW	: in integer range 0 to cFWGlobal;
		   Mult029bFW	: in integer range 0 to cFWGlobal;
		   Mult030bFW	: in integer range 0 to cFWGlobal;
		   Mult031bFW	: in integer range 0 to cFWGlobal;
		   Mult032bFW	: in integer range 0 to cFWGlobal;
		   Mult033bFW	: in integer range 0 to cFWGlobal;
		   Mult034bFW	: in integer range 0 to cFWGlobal;
		   Mult035bFW	: in integer range 0 to cFWGlobal;
		   Mult036bFW	: in integer range 0 to cFWGlobal;
		   Mult037bFW	: in integer range 0 to cFWGlobal;
		   Mult038bFW	: in integer range 0 to cFWGlobal;
		   Mult039bFW	: in integer range 0 to cFWGlobal;
		   Mult040bFW	: in integer range 0 to cFWGlobal;
		   Mult041bFW	: in integer range 0 to cFWGlobal;
		   Mult042bFW	: in integer range 0 to cFWGlobal;
		   Mult043bFW	: in integer range 0 to cFWGlobal;
		   Mult044bFW	: in integer range 0 to cFWGlobal;
		   Mult045bFW	: in integer range 0 to cFWGlobal;
		   Mult046bFW	: in integer range 0 to cFWGlobal;
		   Mult047bFW	: in integer range 0 to cFWGlobal;
		   Mult048bFW	: in integer range 0 to cFWGlobal;
		   Mult049bFW	: in integer range 0 to cFWGlobal;
		   Mult050bFW	: in integer range 0 to cFWGlobal;
		   Mult051bFW	: in integer range 0 to cFWGlobal;
		   Mult052bFW	: in integer range 0 to cFWGlobal;
		   Mult053bFW	: in integer range 0 to cFWGlobal;
		   Mult054bFW	: in integer range 0 to cFWGlobal;
		   Mult055bFW	: in integer range 0 to cFWGlobal;
		   Mult056bFW	: in integer range 0 to cFWGlobal;
		   Mult057bFW	: in integer range 0 to cFWGlobal;
		   Mult058bFW	: in integer range 0 to cFWGlobal;
		   Mult059bFW	: in integer range 0 to cFWGlobal;
		   Mult060bFW	: in integer range 0 to cFWGlobal;
		   Mult061bFW	: in integer range 0 to cFWGlobal;
		   Mult062bFW	: in integer range 0 to cFWGlobal;
		   Mult063bFW	: in integer range 0 to cFWGlobal;
		   Mult064bFW	: in integer range 0 to cFWGlobal;
		   Mult065bFW	: in integer range 0 to cFWGlobal;
		   Mult066bFW	: in integer range 0 to cFWGlobal;
		   Mult067bFW	: in integer range 0 to cFWGlobal;
		   Mult068bFW	: in integer range 0 to cFWGlobal;
		   Mult069bFW	: in integer range 0 to cFWGlobal;
		   Mult070bFW	: in integer range 0 to cFWGlobal;
		   Mult071bFW	: in integer range 0 to cFWGlobal;
		   Mult072bFW	: in integer range 0 to cFWGlobal;
		   Mult073bFW	: in integer range 0 to cFWGlobal;
		   Mult074bFW	: in integer range 0 to cFWGlobal;
		   Mult075bFW	: in integer range 0 to cFWGlobal;
		   Mult076bFW	: in integer range 0 to cFWGlobal;
		   Mult077bFW	: in integer range 0 to cFWGlobal;
		   Mult078bFW	: in integer range 0 to cFWGlobal;
		   Mult079bFW	: in integer range 0 to cFWGlobal;
		   Mult080bFW	: in integer range 0 to cFWGlobal;
		   Mult081bFW	: in integer range 0 to cFWGlobal;
		   Mult082bFW	: in integer range 0 to cFWGlobal;
		   Mult083bFW	: in integer range 0 to cFWGlobal;
		   Mult084bFW	: in integer range 0 to cFWGlobal;
		   Mult085bFW	: in integer range 0 to cFWGlobal;
		   Mult086bFW	: in integer range 0 to cFWGlobal;
		   Mult087bFW	: in integer range 0 to cFWGlobal;
		   Mult088bFW	: in integer range 0 to cFWGlobal;
		   Mult089bFW	: in integer range 0 to cFWGlobal;
		   Mult090bFW	: in integer range 0 to cFWGlobal;
		   Mult091bFW	: in integer range 0 to cFWGlobal;
		   Mult092bFW	: in integer range 0 to cFWGlobal;
		   Mult093bFW	: in integer range 0 to cFWGlobal;
		   Mult094bFW	: in integer range 0 to cFWGlobal;
		   Mult095bFW	: in integer range 0 to cFWGlobal;
		   Mult096bFW	: in integer range 0 to cFWGlobal;
		   Mult097bFW	: in integer range 0 to cFWGlobal;
		   Mult098bFW	: in integer range 0 to cFWGlobal;
		   Mult099bFW	: in integer range 0 to cFWGlobal;
		   Mult100bFW	: in integer range 0 to cFWGlobal;
		   Mult101bFW	: in integer range 0 to cFWGlobal;
		   Mult102bFW	: in integer range 0 to cFWGlobal;
		   Mult103bFW	: in integer range 0 to cFWGlobal;
		   Mult104bFW	: in integer range 0 to cFWGlobal;
		   Mult105bFW	: in integer range 0 to cFWGlobal;
		   Mult106bFW	: in integer range 0 to cFWGlobal;
		   Mult107bFW	: in integer range 0 to cFWGlobal;
		   Mult108bFW	: in integer range 0 to cFWGlobal;
		   Mult109bFW	: in integer range 0 to cFWGlobal;
		   Mult110bFW	: in integer range 0 to cFWGlobal;
		   Mult111bFW	: in integer range 0 to cFWGlobal;
		   Mult112bFW	: in integer range 0 to cFWGlobal;
		   Mult113bFW	: in integer range 0 to cFWGlobal;
		   Mult114bFW	: in integer range 0 to cFWGlobal;
		   Mult115bFW	: in integer range 0 to cFWGlobal;
		   Mult116bFW	: in integer range 0 to cFWGlobal;
		   Mult117bFW	: in integer range 0 to cFWGlobal;
		   Mult118bFW	: in integer range 0 to cFWGlobal;
		   Mult119bFW	: in integer range 0 to cFWGlobal;
		   Mult120bFW	: in integer range 0 to cFWGlobal;
		   Mult121bFW	: in integer range 0 to cFWGlobal;
		   Mult122bFW	: in integer range 0 to cFWGlobal;
		   Mult123bFW	: in integer range 0 to cFWGlobal;
		   Mult124bFW	: in integer range 0 to cFWGlobal;
		   Mult125bFW	: in integer range 0 to cFWGlobal;
		   Mult126bFW	: in integer range 0 to cFWGlobal;
		   Mult127bFW	: in integer range 0 to cFWGlobal;
		   Mult128bFW	: in integer range 0 to cFWGlobal;
		   Mult129bFW	: in integer range 0 to cFWGlobal;
		   Mult130bFW	: in integer range 0 to cFWGlobal;
		   Mult131bFW	: in integer range 0 to cFWGlobal;
		   Mult132bFW	: in integer range 0 to cFWGlobal;
		   Mult133bFW	: in integer range 0 to cFWGlobal;
		   Mult134bFW	: in integer range 0 to cFWGlobal;
		   Mult135bFW	: in integer range 0 to cFWGlobal;
		   Mult136bFW	: in integer range 0 to cFWGlobal;
		   Mult137bFW	: in integer range 0 to cFWGlobal;
		   Mult138bFW	: in integer range 0 to cFWGlobal;
		   Mult139bFW	: in integer range 0 to cFWGlobal;
		   Mult140bFW	: in integer range 0 to cFWGlobal;
		   Mult141bFW	: in integer range 0 to cFWGlobal;
		   Mult142bFW	: in integer range 0 to cFWGlobal;
		   Mult143bFW	: in integer range 0 to cFWGlobal;
		   Mult144bFW	: in integer range 0 to cFWGlobal;
		   Mult145bFW	: in integer range 0 to cFWGlobal;
		   Mult146bFW	: in integer range 0 to cFWGlobal;
		   Mult147bFW	: in integer range 0 to cFWGlobal;
		   Mult148bFW	: in integer range 0 to cFWGlobal;
		   Mult149bFW	: in integer range 0 to cFWGlobal;
		   Mult150bFW	: in integer range 0 to cFWGlobal
		);
		   
		   
end FIR_Example;

architecture Behavioral of FIR_Example is
	-- Coefficients 
    constant Coeff000 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111101100011111001000100110";
    constant Coeff001 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111110111101011101010011111000";
    constant Coeff002 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111101001011010101001011001";
    constant Coeff003 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000100111100001000101001011";
    constant Coeff004 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000101010001110101010011011";
    constant Coeff005 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111111010100100011010111100";
    constant Coeff006 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111011000110111100101101100";
    constant Coeff007 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111101010001101100000001010";
    constant Coeff008 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000010100111001000001011000";
    constant Coeff009 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000100011010011101110100111";
    constant Coeff010 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000011001011010011101000";
    constant Coeff011 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111011101110101100110000011";
    constant Coeff012 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111100110100100001000001001";
    constant Coeff013 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000010100010101101010010010";
    constant Coeff014 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000100111111110011100011011";
    constant Coeff015 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000010100000011001101100";
    constant Coeff016 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111010110001001000101110101";
    constant Coeff017 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111100011101011110101110000";
    constant Coeff018 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000011100000110010010110100";
    constant Coeff019 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000110000001100110001110100";
    constant Coeff020 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111111111101001000000111000";
    constant Coeff021 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111001011011010000011001010";
    constant Coeff022 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111011110110101111010101010";
    constant Coeff023 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000100011110101110011111011";
    constant Coeff024 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000111011001101101111001111";
    constant Coeff025 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111111111011101011010001000";
    constant Coeff026 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111110111111001111111110101011";
    constant Coeff027 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111010110011101000010010101";
    constant Coeff028 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000101011010111101011101111";
    constant Coeff029 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000001001001010010001111010110";
    constant Coeff030 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000000011001110001101010";
    constant Coeff031 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111110110000110011010001100000";
    constant Coeff032 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111001100011110110011010011";
    constant Coeff033 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000110100100010101111000101";
    constant Coeff034 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000001011001100000100110100001";
    constant Coeff035 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000000101101000000110011";
    constant Coeff036 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111110011111101010111100110010";
    constant Coeff037 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111000001010110110111000010";
    constant Coeff038 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000001000000000000001000110110";
    constant Coeff039 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000001101101000001001100011010";
    constant Coeff040 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000000101110111110000010";
    constant Coeff041 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111110001010000101000111001010";
    constant Coeff042 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111110110011001101111000101000";
    constant Coeff043 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000001001110111010000101110010";
    constant Coeff044 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000010000110101001101110010101";
    constant Coeff045 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000000110000100100101001";
    constant Coeff046 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111101101101001101110111000110";
    constant Coeff047 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111110100000010000101000001001";
    constant Coeff048 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000001100011000100111110011011";
    constant Coeff049 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000010101001011001100101100100";
    constant Coeff050 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000000110001011110100111";
    constant Coeff051 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111101000101100101011000000100";
    constant Coeff052 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111110000101111010010101011011";
    constant Coeff053 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000001111111001110110100100001";
    constant Coeff054 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000011011010110110110010010000";
    constant Coeff055 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000001000001101011010110";
    constant Coeff056 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111100001011010101001101010011";
    constant Coeff057 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111101011110001011000111001110";
    constant Coeff058 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000010101010011001100001001100";
    constant Coeff059 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000100101000110001001011111000";
    constant Coeff060 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000001010101000000001110";
    constant Coeff061 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111010101010001000000111111110";
    constant Coeff062 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111100011001111111100010001101";
    constant Coeff063 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000011110111111100110111001001";
    constant Coeff064 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000110111001110011110111101111";
    constant Coeff065 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000001010110001010101111";
    constant Coeff066 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111110111100001001010000000110010";
    constant Coeff067 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111010000100000110010111111001";
    constant Coeff068 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000110110001000011111011110110";
    constant Coeff069 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000001100110101101111001100110100";
    constant Coeff070 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000001010000110111011000";
    constant Coeff071 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111101100101011111110101001100010";
    constant Coeff072 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111110000000010110110001100010001";
    constant Coeff073 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000010111111010100101001101111100";
    constant Coeff074 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000001001101011111011011001010000100";
    constant Coeff075 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000001100110011010110110011000111101";
    constant Coeff076 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000001001101011111011011001010000100";
    constant Coeff077 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000010111111010100101001101111100";
    constant Coeff078 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111110000000010110110001100010001";
    constant Coeff079 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111101100101011111110101001100010";
    constant Coeff080 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000001010000110111011000";
    constant Coeff081 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000001100110101101111001100110100";
    constant Coeff082 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000110110001000011111011110110";
    constant Coeff083 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111010000100000110010111111001";
    constant Coeff084 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111110111100001001010000000110010";
    constant Coeff085 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000001010110001010101111";
    constant Coeff086 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000110111001110011110111101111";
    constant Coeff087 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000011110111111100110111001001";
    constant Coeff088 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111100011001111111100010001101";
    constant Coeff089 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111010101010001000000111111110";
    constant Coeff090 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000001010101000000001110";
    constant Coeff091 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000100101000110001001011111000";
    constant Coeff092 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000010101010011001100001001100";
    constant Coeff093 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111101011110001011000111001110";
    constant Coeff094 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111100001011010101001101010011";
    constant Coeff095 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000001000001101011010110";
    constant Coeff096 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000011011010110110110010010000";
    constant Coeff097 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000001111111001110110100100001";
    constant Coeff098 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111110000101111010010101011011";
    constant Coeff099 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111101000101100101011000000100";
    constant Coeff100 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000000110001011110100111";
    constant Coeff101 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000010101001011001100101100100";
    constant Coeff102 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000001100011000100111110011011";
    constant Coeff103 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111110100000010000101000001001";
    constant Coeff104 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111101101101001101110111000110";
    constant Coeff105 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000000110000100100101001";
    constant Coeff106 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000010000110101001101110010101";
    constant Coeff107 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000001001110111010000101110010";
    constant Coeff108 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111110110011001101111000101000";
    constant Coeff109 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111110001010000101000111001010";
    constant Coeff110 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000000101110111110000010";
    constant Coeff111 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000001101101000001001100011010";
    constant Coeff112 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000001000000000000001000110110";
    constant Coeff113 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111000001010110110111000010";
    constant Coeff114 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111110011111101010111100110010";
    constant Coeff115 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000000101101000000110011";
    constant Coeff116 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000001011001100000100110100001";
    constant Coeff117 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000110100100010101111000101";
    constant Coeff118 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111001100011110110011010011";
    constant Coeff119 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111110110000110011010001100000";
    constant Coeff120 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000000011001110001101010";
    constant Coeff121 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000001001001010010001111010110";
    constant Coeff122 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000101011010111101011101111";
    constant Coeff123 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111010110011101000010010101";
    constant Coeff124 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111110111111001111111110101011";
    constant Coeff125 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111111111011101011010001000";
    constant Coeff126 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000111011001101101111001111";
    constant Coeff127 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000100011110101110011111011";
    constant Coeff128 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111011110110101111010101010";
    constant Coeff129 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111001011011010000011001010";
    constant Coeff130 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111111111101001000000111000";
    constant Coeff131 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000110000001100110001110100";
    constant Coeff132 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000011100000110010010110100";
    constant Coeff133 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111100011101011110101110000";
    constant Coeff134 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111010110001001000101110101";
    constant Coeff135 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000010100000011001101100";
    constant Coeff136 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000100111111110011100011011";
    constant Coeff137 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000010100010101101010010010";
    constant Coeff138 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111100110100100001000001001";
    constant Coeff139 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111011101110101100110000011";
    constant Coeff140 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000000011001011010011101000";
    constant Coeff141 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000100011010011101110100111";
    constant Coeff142 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000010100111001000001011000";
    constant Coeff143 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111101010001101100000001010";
    constant Coeff144 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111011000110111100101101100";
    constant Coeff145 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111111010100100011010111100";
    constant Coeff146 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000101010001110101010011011";
    constant Coeff147 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "0000000000000000000000000000000000000000100111100001000101001011";
    constant Coeff148 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111101001011010101001011001";
    constant Coeff149 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111110111101011101010011111000";
    constant Coeff150 : Signed (cIWGlobal+cFWGlobal-1 downto 0) := "1111111111111111111111111111111111111111101100011111001000100110";
	
	-- input delay line
	signal X000	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X001	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X002	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X003	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X004	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X005	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X006	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X007	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X008	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X009	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X010	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X011	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X012	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X013	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X014	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X015	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X016	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X017	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X018	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X019	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X020	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X021	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X022	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X023	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X024	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X025	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X026	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X027	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X028	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X029	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X030	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X031	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X032	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X033	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X034	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X035	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X036	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X037	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X038	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X039	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X040	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X041	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X042	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X043	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X044	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X045	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X046	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X047	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X048	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X049	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X050	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X051	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X052	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X053	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X054	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X055	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X056	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X057	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X058	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X059	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X060	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X061	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X062	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X063	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X064	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X065	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X066	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X067	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X068	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X069	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X070	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X071	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X072	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X073	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X074	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X075	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X076	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X077	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X078	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X079	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X080	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X081	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X082	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X083	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X084	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X085	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X086	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X087	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X088	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X089	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X090	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X091	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X092	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X093	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X094	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X095	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X096	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X097	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X098	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X099	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X100	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X101	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X102	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X103	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X104	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X105	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X106	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X107	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X108	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X109	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X110	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X111	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X112	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X113	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X114	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X115	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X116	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X117	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X118	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X119	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X120	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X121	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X122	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X123	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X124	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X125	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X126	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X127	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X128	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X129	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X130	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X131	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X132	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X133	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X134	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X135	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X136	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X137	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X138	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X139	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X140	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X141	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X142	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X143	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X144	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X145	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X146	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X147	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X148	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X149	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal X150	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');


	constant Y000	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y001	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y002	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y003	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y004	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y005	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y006	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y007	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y008	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y009	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y010	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y011	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y012	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y013	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y014	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y015	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y016	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y017	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y018	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y019	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y020	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y021	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y022	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y023	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y024	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y025	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y026	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y027	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y028	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y029	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y030	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y031	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y032	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y033	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y034	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y035	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y036	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y037	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y038	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y039	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y040	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y041	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y042	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y043	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y044	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y045	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y046	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y047	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y048	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y049	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y050	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y051	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y052	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y053	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y054	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y055	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y056	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y057	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y058	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y059	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y060	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y061	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y062	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y063	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y064	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y065	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y066	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y067	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y068	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y069	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y070	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y071	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y072	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y073	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y074	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y075	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y076	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y077	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y078	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y079	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y080	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y081	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y082	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y083	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y084	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y085	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y086	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y087	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y088	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y089	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y090	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y091	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y092	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y093	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y094	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y095	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y096	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y097	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y098	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y099	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y100	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y101	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y102	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y103	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y104	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y105	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y106	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y107	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y108	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y109	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y110	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y111	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y112	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y113	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y114	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y115	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y116	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y117	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y118	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y119	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y120	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y121	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y122	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y123	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y124	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y125	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y126	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y127	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y128	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y129	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y130	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y131	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y132	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y133	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y134	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y135	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y136	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y137	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y138	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y139	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y140	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y141	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y142	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y143	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y144	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y145	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y146	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y147	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y148	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y149	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal Y150	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	
	--Multiply Output
	signal MultOut000  	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut001  	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut002  	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut003  	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut004  	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut005  	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut006  	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut007  	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut008  	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut009  	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut010 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut011 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut012 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut013 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut014 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut015 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut016 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut017 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut018 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut019 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut020 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut021 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut022 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut023 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut024 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut025 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut026 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut027 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut028 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut029 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut030 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut031 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut032 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut033 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut034 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut035 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut036 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut037 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut038 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut039 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut040 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut041 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut042 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut043 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut044 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut045 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut046 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut047 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut048 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut049 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut050 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut051 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut052 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut053 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut054 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut055 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut056 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut057 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut058 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut059 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut060 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut061 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut062 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut063 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut064 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut065 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut066 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut067 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut068 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut069 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut070 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut071 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut072 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut073 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut074 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut075 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut076 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut077 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut078 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut079 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut080 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut081 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut082 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut083 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut084 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut085 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut086 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut087 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut088 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut089 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut090 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut091 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut092 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut093 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut094 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut095 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut096 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut097 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut098 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut099 	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut100	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut101	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut102	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut103	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut104	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut105	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut106	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut107	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut108	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut109	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut110	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut111	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut112	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut113	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut114	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut115	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut116	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut117	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut118	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut119	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut120	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut121	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut122	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut123	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut124	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut125	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut126	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut127	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut128	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut129	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut130	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut131	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut132	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut133	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut134	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut135	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut136	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut137	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut138	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut139	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut140	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut141	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut142	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut143	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut144	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut145	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut146	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut147	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut148	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut149	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');
	signal MultOut150	: Signed (cIWGlobal+cFWGlobal-1 downto 0) := (others => '0');

	component WC_Mult is
		Generic(
			cIWGlobal		: integer := 32; --Input Integer part Width
			cFWGlobal		: integer := 32 --Input Fractional part Width
			);
		Port ( 
			I1 : in signed (cIWGlobal+cFWGlobal-1 downto 0);
			I2 : in signed (cIWGlobal+cFWGlobal-1 downto 0);
			O : out signed (cIWGlobal+cFWGlobal-1 downto 0);
	
			-- Widths for the Width Adapters
	
			In1IW	: in integer range 0 to cIWGlobal; --Output Integer part Width
			In1FW	: in integer range 0 to cFWGlobal; --Output Fractional part Width
			In2IW	: in integer range 0 to cIWGlobal; --Output Integer part Width
			In2FW	: in integer range 0 to cFWGlobal --Output Fractional part Width
	
			);
	end component WC_Mult;
	
	component WC_AddSub is
		Generic(
			cIWGlobal		: integer := 32; --Input Integer part Width
			cFWGlobal		: integer := 32; --Input Fractional part Width
			cAddSubSel		: boolean := true --Add/Subtract Select
			);
		Port ( 
			I1 : in signed (cIWGlobal+cFWGlobal-1 downto 0);
			I2 : in signed (cIWGlobal+cFWGlobal-1 downto 0);
			O : out signed (cIWGlobal+cFWGlobal-1 downto 0);
	
			-- Widths for the Width Adapters
	
			In1IW	: in integer range 0 to cIWGlobal; --Output Integer part Width
			In1FW	: in integer range 0 to cFWGlobal; --Output Fractional part Width
			In2IW	: in integer range 0 to cIWGlobal; --Output Integer part Width
			In2FW	: in integer range 0 to cFWGlobal --Output Fractional part Width
	
			);
	end component WC_AddSub;
	
	
begin
	
	-- input delay line process structure
	X000	<=	X;

	process (Clk)
	begin
	if (Clk'event and Clk = '1') then
		if Rst = '0' then
		--	X000 <= (others => '0'); X0 is alias to X
			X001 <= (others => '0');
			X002 <= (others => '0');
			X003 <= (others => '0');
			X004 <= (others => '0');
			X005 <= (others => '0');
			X006 <= (others => '0');
			X007 <= (others => '0');
			X008 <= (others => '0');
			X009 <= (others => '0');
			X010 <= (others => '0');
			X011 <= (others => '0');
			X012 <= (others => '0');
			X013 <= (others => '0');
			X014 <= (others => '0');
			X015 <= (others => '0');
			X016 <= (others => '0');
			X017 <= (others => '0');
			X018 <= (others => '0');
			X019 <= (others => '0');
			X020 <= (others => '0');
			X021 <= (others => '0');
			X022 <= (others => '0');
			X023 <= (others => '0');
			X024 <= (others => '0');
			X025 <= (others => '0');
			X026 <= (others => '0');
			X027 <= (others => '0');
			X028 <= (others => '0');
			X029 <= (others => '0');
			X030 <= (others => '0');
			X031 <= (others => '0');
			X032 <= (others => '0');
			X033 <= (others => '0');
			X034 <= (others => '0');
			X035 <= (others => '0');
			X036 <= (others => '0');
			X037 <= (others => '0');
			X038 <= (others => '0');
			X039 <= (others => '0');
			X040 <= (others => '0');
			X041 <= (others => '0');
			X042 <= (others => '0');
			X043 <= (others => '0');
			X044 <= (others => '0');
			X045 <= (others => '0');
			X046 <= (others => '0');
			X047 <= (others => '0');
			X048 <= (others => '0');
			X049 <= (others => '0');
			X050 <= (others => '0');
			X051 <= (others => '0');
			X052 <= (others => '0');
			X053 <= (others => '0');
			X054 <= (others => '0');
			X055 <= (others => '0');
			X056 <= (others => '0');
			X057 <= (others => '0');
			X058 <= (others => '0');
			X059 <= (others => '0');
			X060 <= (others => '0');
			X061 <= (others => '0');
			X062 <= (others => '0');
			X063 <= (others => '0');
			X064 <= (others => '0');
			X065 <= (others => '0');
			X066 <= (others => '0');
			X067 <= (others => '0');
			X068 <= (others => '0');
			X069 <= (others => '0');
			X070 <= (others => '0');
			X071 <= (others => '0');
			X072 <= (others => '0');
			X073 <= (others => '0');
			X074 <= (others => '0');
			X075 <= (others => '0');
			X076 <= (others => '0');
			X077 <= (others => '0');
			X078 <= (others => '0');
			X079 <= (others => '0');
			X080 <= (others => '0');
			X081 <= (others => '0');
			X082 <= (others => '0');
			X083 <= (others => '0');
			X084 <= (others => '0');
			X085 <= (others => '0');
			X086 <= (others => '0');
			X087 <= (others => '0');
			X088 <= (others => '0');
			X089 <= (others => '0');
			X090 <= (others => '0');
			X091 <= (others => '0');
			X092 <= (others => '0');
			X093 <= (others => '0');
			X094 <= (others => '0');
			X095 <= (others => '0');
			X096 <= (others => '0');
			X097 <= (others => '0');
			X098 <= (others => '0');
			X099 <= (others => '0');
			X100 <= (others => '0');
			X101 <= (others => '0');
			X102 <= (others => '0');
			X103 <= (others => '0');
			X104 <= (others => '0');
			X105 <= (others => '0');
			X106 <= (others => '0');
			X107 <= (others => '0');
			X108 <= (others => '0');
			X109 <= (others => '0');
			X110 <= (others => '0');
			X111 <= (others => '0');
			X112 <= (others => '0');
			X113 <= (others => '0');
			X114 <= (others => '0');
			X115 <= (others => '0');
			X116 <= (others => '0');
			X117 <= (others => '0');
			X118 <= (others => '0');
			X119 <= (others => '0');
			X120 <= (others => '0');
			X121 <= (others => '0');
			X122 <= (others => '0');
			X123 <= (others => '0');
			X124 <= (others => '0');
			X125 <= (others => '0');
			X126 <= (others => '0');
			X127 <= (others => '0');
			X128 <= (others => '0');
			X129 <= (others => '0');
			X130 <= (others => '0');
			X131 <= (others => '0');
			X132 <= (others => '0');
			X133 <= (others => '0');
			X134 <= (others => '0');
			X135 <= (others => '0');
			X136 <= (others => '0');
			X137 <= (others => '0');
			X138 <= (others => '0');
			X139 <= (others => '0');
			X140 <= (others => '0');
			X141 <= (others => '0');
			X142 <= (others => '0');
			X143 <= (others => '0');
			X144 <= (others => '0');
			X145 <= (others => '0');
			X146 <= (others => '0');
			X147 <= (others => '0');
			X148 <= (others => '0');
			X149 <= (others => '0');
			X150 <= (others => '0');
		else
			--X000 <= X;
			X001 <= X000;
			X002 <= X001;
			X003 <= X002;
			X004 <= X003;
			X005 <= X004;
			X006 <= X005;
			X007 <= X006;
			X008 <= X007;
			X009 <= X008;
			X010 <= X009;
			X011 <= X010;
			X012 <= X011;
			X013 <= X012;
			X014 <= X013;
			X015 <= X014;
			X016 <= X015;
			X017 <= X016;
			X018 <= X017;
			X019 <= X018;
			X020 <= X019;
			X021 <= X020;
			X022 <= X021;
			X023 <= X022;
			X024 <= X023;
			X025 <= X024;
			X026 <= X025;
			X027 <= X026;
			X028 <= X027;
			X029 <= X028;
			X030 <= X029;
			X031 <= X030;
			X032 <= X031;
			X033 <= X032;
			X034 <= X033;
			X035 <= X034;
			X036 <= X035;
			X037 <= X036;
			X038 <= X037;
			X039 <= X038;
			X040 <= X039;
			X041 <= X040;
			X042 <= X041;
			X043 <= X042;
			X044 <= X043;
			X045 <= X044;
			X046 <= X045;
			X047 <= X046;
			X048 <= X047;
			X049 <= X048;
			X050 <= X049;
			X051 <= X050;
			X052 <= X051;
			X053 <= X052;
			X054 <= X053;
			X055 <= X054;
			X056 <= X055;
			X057 <= X056;
			X058 <= X057;
			X059 <= X058;
			X060 <= X059;
			X061 <= X060;
			X062 <= X061;
			X063 <= X062;
			X064 <= X063;
			X065 <= X064;
			X066 <= X065;
			X067 <= X066;
			X068 <= X067;
			X069 <= X068;
			X070 <= X069;
			X071 <= X070;
			X072 <= X071;
			X073 <= X072;
			X074 <= X073;
			X075 <= X074;
			X076 <= X075;
			X077 <= X076;
			X078 <= X077;
			X079 <= X078;
			X080 <= X079;
			X081 <= X080;
			X082 <= X081;
			X083 <= X082;
			X084 <= X083;
			X085 <= X084;
			X086 <= X085;
			X087 <= X086;
			X088 <= X087;
			X089 <= X088;
			X090 <= X089;
			X091 <= X090;
			X092 <= X091;
			X093 <= X092;
			X094 <= X093;
			X095 <= X094;
			X096 <= X095;
			X097 <= X096;
			X098 <= X097;
			X099 <= X098;
			X100 <= X099;
			X101 <= X100;
			X102 <= X101;
			X103 <= X102;
			X104 <= X103;
			X105 <= X104;
			X106 <= X105;
			X107 <= X106;
			X108 <= X107;
			X109 <= X108;
			X110 <= X109;
			X111 <= X110;
			X112 <= X111;
			X113 <= X112;
			X114 <= X113;
			X115 <= X114;
			X116 <= X115;
			X117 <= X116;
			X118 <= X117;
			X119 <= X118;
			X120 <= X119;
			X121 <= X120;
			X122 <= X121;
			X123 <= X122;
			X124 <= X123;
			X125 <= X124;
			X126 <= X125;
			X127 <= X126;
			X128 <= X127;
			X129 <= X128;
			X130 <= X129;
			X131 <= X130;
			X132 <= X131;
			X133 <= X132;
			X134 <= X133;
			X135 <= X134;
			X136 <= X135;
			X137 <= X136;
			X138 <= X137;
			X139 <= X138;
			X140 <= X139;
			X141 <= X140;
			X142 <= X141;
			X143 <= X142;
			X144 <= X143;
			X145 <= X144;
			X146 <= X145;
			X147 <= X146;
			X148 <= X147;
			X149 <= X148;
			X150 <= X149;
		end if;
	end if;
	end process;

	-- Multipliers
	WC_Mult000:	WC_Mult port map (I1 => X000, I2 => Coeff000, O => MultOut000, In1IW => Mult000aIW, In1FW => Mult000aFW, In2IW => Mult000bIW, In2FW => Mult000bFW);
	WC_Mult001:	WC_Mult port map (I1 => X001, I2 => Coeff001, O => MultOut001, In1IW => Mult001aIW, In1FW => Mult001aFW, In2IW => Mult001bIW, In2FW => Mult001bFW);
	WC_Mult002:	WC_Mult port map (I1 => X002, I2 => Coeff002, O => MultOut002, In1IW => Mult002aIW, In1FW => Mult002aFW, In2IW => Mult002bIW, In2FW => Mult002bFW);
	WC_Mult003:	WC_Mult port map (I1 => X003, I2 => Coeff003, O => MultOut003, In1IW => Mult003aIW, In1FW => Mult003aFW, In2IW => Mult003bIW, In2FW => Mult003bFW);
	WC_Mult004:	WC_Mult port map (I1 => X004, I2 => Coeff004, O => MultOut004, In1IW => Mult004aIW, In1FW => Mult004aFW, In2IW => Mult004bIW, In2FW => Mult004bFW);
	WC_Mult005:	WC_Mult port map (I1 => X005, I2 => Coeff005, O => MultOut005, In1IW => Mult005aIW, In1FW => Mult005aFW, In2IW => Mult005bIW, In2FW => Mult005bFW);
	WC_Mult006:	WC_Mult port map (I1 => X006, I2 => Coeff006, O => MultOut006, In1IW => Mult006aIW, In1FW => Mult006aFW, In2IW => Mult006bIW, In2FW => Mult006bFW);
	WC_Mult007:	WC_Mult port map (I1 => X007, I2 => Coeff007, O => MultOut007, In1IW => Mult007aIW, In1FW => Mult007aFW, In2IW => Mult007bIW, In2FW => Mult007bFW);
	WC_Mult008:	WC_Mult port map (I1 => X008, I2 => Coeff008, O => MultOut008, In1IW => Mult008aIW, In1FW => Mult008aFW, In2IW => Mult008bIW, In2FW => Mult008bFW);
	WC_Mult009:	WC_Mult port map (I1 => X009, I2 => Coeff009, O => MultOut009, In1IW => Mult009aIW, In1FW => Mult009aFW, In2IW => Mult009bIW, In2FW => Mult009bFW);
	WC_Mult010:	WC_Mult port map (I1 => X010, I2 => Coeff010, O => MultOut010, In1IW => Mult010aIW, In1FW => Mult010aFW, In2IW => Mult010bIW, In2FW => Mult010bFW);
	WC_Mult011:	WC_Mult port map (I1 => X011, I2 => Coeff011, O => MultOut011, In1IW => Mult011aIW, In1FW => Mult011aFW, In2IW => Mult011bIW, In2FW => Mult011bFW);
	WC_Mult012:	WC_Mult port map (I1 => X012, I2 => Coeff012, O => MultOut012, In1IW => Mult012aIW, In1FW => Mult012aFW, In2IW => Mult012bIW, In2FW => Mult012bFW);
	WC_Mult013:	WC_Mult port map (I1 => X013, I2 => Coeff013, O => MultOut013, In1IW => Mult013aIW, In1FW => Mult013aFW, In2IW => Mult013bIW, In2FW => Mult013bFW);
	WC_Mult014:	WC_Mult port map (I1 => X014, I2 => Coeff014, O => MultOut014, In1IW => Mult014aIW, In1FW => Mult014aFW, In2IW => Mult014bIW, In2FW => Mult014bFW);
	WC_Mult015:	WC_Mult port map (I1 => X015, I2 => Coeff015, O => MultOut015, In1IW => Mult015aIW, In1FW => Mult015aFW, In2IW => Mult015bIW, In2FW => Mult015bFW);
	WC_Mult016:	WC_Mult port map (I1 => X016, I2 => Coeff016, O => MultOut016, In1IW => Mult016aIW, In1FW => Mult016aFW, In2IW => Mult016bIW, In2FW => Mult016bFW);
	WC_Mult017:	WC_Mult port map (I1 => X017, I2 => Coeff017, O => MultOut017, In1IW => Mult017aIW, In1FW => Mult017aFW, In2IW => Mult017bIW, In2FW => Mult017bFW);
	WC_Mult018:	WC_Mult port map (I1 => X018, I2 => Coeff018, O => MultOut018, In1IW => Mult018aIW, In1FW => Mult018aFW, In2IW => Mult018bIW, In2FW => Mult018bFW);
	WC_Mult019:	WC_Mult port map (I1 => X019, I2 => Coeff019, O => MultOut019, In1IW => Mult019aIW, In1FW => Mult019aFW, In2IW => Mult019bIW, In2FW => Mult019bFW);
	WC_Mult020:	WC_Mult port map (I1 => X020, I2 => Coeff020, O => MultOut020, In1IW => Mult020aIW, In1FW => Mult020aFW, In2IW => Mult020bIW, In2FW => Mult020bFW);
	WC_Mult021:	WC_Mult port map (I1 => X021, I2 => Coeff021, O => MultOut021, In1IW => Mult021aIW, In1FW => Mult021aFW, In2IW => Mult021bIW, In2FW => Mult021bFW);
	WC_Mult022:	WC_Mult port map (I1 => X022, I2 => Coeff022, O => MultOut022, In1IW => Mult022aIW, In1FW => Mult022aFW, In2IW => Mult022bIW, In2FW => Mult022bFW);
	WC_Mult023:	WC_Mult port map (I1 => X023, I2 => Coeff023, O => MultOut023, In1IW => Mult023aIW, In1FW => Mult023aFW, In2IW => Mult023bIW, In2FW => Mult023bFW);
	WC_Mult024:	WC_Mult port map (I1 => X024, I2 => Coeff024, O => MultOut024, In1IW => Mult024aIW, In1FW => Mult024aFW, In2IW => Mult024bIW, In2FW => Mult024bFW);
	WC_Mult025:	WC_Mult port map (I1 => X025, I2 => Coeff025, O => MultOut025, In1IW => Mult025aIW, In1FW => Mult025aFW, In2IW => Mult025bIW, In2FW => Mult025bFW);
	WC_Mult026:	WC_Mult port map (I1 => X026, I2 => Coeff026, O => MultOut026, In1IW => Mult026aIW, In1FW => Mult026aFW, In2IW => Mult026bIW, In2FW => Mult026bFW);
	WC_Mult027:	WC_Mult port map (I1 => X027, I2 => Coeff027, O => MultOut027, In1IW => Mult027aIW, In1FW => Mult027aFW, In2IW => Mult027bIW, In2FW => Mult027bFW);
	WC_Mult028:	WC_Mult port map (I1 => X028, I2 => Coeff028, O => MultOut028, In1IW => Mult028aIW, In1FW => Mult028aFW, In2IW => Mult028bIW, In2FW => Mult028bFW);
	WC_Mult029:	WC_Mult port map (I1 => X029, I2 => Coeff029, O => MultOut029, In1IW => Mult029aIW, In1FW => Mult029aFW, In2IW => Mult029bIW, In2FW => Mult029bFW);
	WC_Mult030:	WC_Mult port map (I1 => X030, I2 => Coeff030, O => MultOut030, In1IW => Mult030aIW, In1FW => Mult030aFW, In2IW => Mult030bIW, In2FW => Mult030bFW);
	WC_Mult031:	WC_Mult port map (I1 => X031, I2 => Coeff031, O => MultOut031, In1IW => Mult031aIW, In1FW => Mult031aFW, In2IW => Mult031bIW, In2FW => Mult031bFW);
	WC_Mult032:	WC_Mult port map (I1 => X032, I2 => Coeff032, O => MultOut032, In1IW => Mult032aIW, In1FW => Mult032aFW, In2IW => Mult032bIW, In2FW => Mult032bFW);
	WC_Mult033:	WC_Mult port map (I1 => X033, I2 => Coeff033, O => MultOut033, In1IW => Mult033aIW, In1FW => Mult033aFW, In2IW => Mult033bIW, In2FW => Mult033bFW);
	WC_Mult034:	WC_Mult port map (I1 => X034, I2 => Coeff034, O => MultOut034, In1IW => Mult034aIW, In1FW => Mult034aFW, In2IW => Mult034bIW, In2FW => Mult034bFW);
	WC_Mult035:	WC_Mult port map (I1 => X035, I2 => Coeff035, O => MultOut035, In1IW => Mult035aIW, In1FW => Mult035aFW, In2IW => Mult035bIW, In2FW => Mult035bFW);
	WC_Mult036:	WC_Mult port map (I1 => X036, I2 => Coeff036, O => MultOut036, In1IW => Mult036aIW, In1FW => Mult036aFW, In2IW => Mult036bIW, In2FW => Mult036bFW);
	WC_Mult037:	WC_Mult port map (I1 => X037, I2 => Coeff037, O => MultOut037, In1IW => Mult037aIW, In1FW => Mult037aFW, In2IW => Mult037bIW, In2FW => Mult037bFW);
	WC_Mult038:	WC_Mult port map (I1 => X038, I2 => Coeff038, O => MultOut038, In1IW => Mult038aIW, In1FW => Mult038aFW, In2IW => Mult038bIW, In2FW => Mult038bFW);
	WC_Mult039:	WC_Mult port map (I1 => X039, I2 => Coeff039, O => MultOut039, In1IW => Mult039aIW, In1FW => Mult039aFW, In2IW => Mult039bIW, In2FW => Mult039bFW);
	WC_Mult040:	WC_Mult port map (I1 => X040, I2 => Coeff040, O => MultOut040, In1IW => Mult040aIW, In1FW => Mult040aFW, In2IW => Mult040bIW, In2FW => Mult040bFW);
	WC_Mult041:	WC_Mult port map (I1 => X041, I2 => Coeff041, O => MultOut041, In1IW => Mult041aIW, In1FW => Mult041aFW, In2IW => Mult041bIW, In2FW => Mult041bFW);
	WC_Mult042:	WC_Mult port map (I1 => X042, I2 => Coeff042, O => MultOut042, In1IW => Mult042aIW, In1FW => Mult042aFW, In2IW => Mult042bIW, In2FW => Mult042bFW);
	WC_Mult043:	WC_Mult port map (I1 => X043, I2 => Coeff043, O => MultOut043, In1IW => Mult043aIW, In1FW => Mult043aFW, In2IW => Mult043bIW, In2FW => Mult043bFW);
	WC_Mult044:	WC_Mult port map (I1 => X044, I2 => Coeff044, O => MultOut044, In1IW => Mult044aIW, In1FW => Mult044aFW, In2IW => Mult044bIW, In2FW => Mult044bFW);
	WC_Mult045:	WC_Mult port map (I1 => X045, I2 => Coeff045, O => MultOut045, In1IW => Mult045aIW, In1FW => Mult045aFW, In2IW => Mult045bIW, In2FW => Mult045bFW);
	WC_Mult046:	WC_Mult port map (I1 => X046, I2 => Coeff046, O => MultOut046, In1IW => Mult046aIW, In1FW => Mult046aFW, In2IW => Mult046bIW, In2FW => Mult046bFW);
	WC_Mult047:	WC_Mult port map (I1 => X047, I2 => Coeff047, O => MultOut047, In1IW => Mult047aIW, In1FW => Mult047aFW, In2IW => Mult047bIW, In2FW => Mult047bFW);
	WC_Mult048:	WC_Mult port map (I1 => X048, I2 => Coeff048, O => MultOut048, In1IW => Mult048aIW, In1FW => Mult048aFW, In2IW => Mult048bIW, In2FW => Mult048bFW);
	WC_Mult049:	WC_Mult port map (I1 => X049, I2 => Coeff049, O => MultOut049, In1IW => Mult049aIW, In1FW => Mult049aFW, In2IW => Mult049bIW, In2FW => Mult049bFW);
	WC_Mult050:	WC_Mult port map (I1 => X050, I2 => Coeff050, O => MultOut050, In1IW => Mult050aIW, In1FW => Mult050aFW, In2IW => Mult050bIW, In2FW => Mult050bFW);
	WC_Mult051:	WC_Mult port map (I1 => X051, I2 => Coeff051, O => MultOut051, In1IW => Mult051aIW, In1FW => Mult051aFW, In2IW => Mult051bIW, In2FW => Mult051bFW);
	WC_Mult052:	WC_Mult port map (I1 => X052, I2 => Coeff052, O => MultOut052, In1IW => Mult052aIW, In1FW => Mult052aFW, In2IW => Mult052bIW, In2FW => Mult052bFW);
	WC_Mult053:	WC_Mult port map (I1 => X053, I2 => Coeff053, O => MultOut053, In1IW => Mult053aIW, In1FW => Mult053aFW, In2IW => Mult053bIW, In2FW => Mult053bFW);
	WC_Mult054:	WC_Mult port map (I1 => X054, I2 => Coeff054, O => MultOut054, In1IW => Mult054aIW, In1FW => Mult054aFW, In2IW => Mult054bIW, In2FW => Mult054bFW);
	WC_Mult055:	WC_Mult port map (I1 => X055, I2 => Coeff055, O => MultOut055, In1IW => Mult055aIW, In1FW => Mult055aFW, In2IW => Mult055bIW, In2FW => Mult055bFW);
	WC_Mult056:	WC_Mult port map (I1 => X056, I2 => Coeff056, O => MultOut056, In1IW => Mult056aIW, In1FW => Mult056aFW, In2IW => Mult056bIW, In2FW => Mult056bFW);
	WC_Mult057:	WC_Mult port map (I1 => X057, I2 => Coeff057, O => MultOut057, In1IW => Mult057aIW, In1FW => Mult057aFW, In2IW => Mult057bIW, In2FW => Mult057bFW);
	WC_Mult058:	WC_Mult port map (I1 => X058, I2 => Coeff058, O => MultOut058, In1IW => Mult058aIW, In1FW => Mult058aFW, In2IW => Mult058bIW, In2FW => Mult058bFW);
	WC_Mult059:	WC_Mult port map (I1 => X059, I2 => Coeff059, O => MultOut059, In1IW => Mult059aIW, In1FW => Mult059aFW, In2IW => Mult059bIW, In2FW => Mult059bFW);
	WC_Mult060:	WC_Mult port map (I1 => X060, I2 => Coeff060, O => MultOut060, In1IW => Mult060aIW, In1FW => Mult060aFW, In2IW => Mult060bIW, In2FW => Mult060bFW);
	WC_Mult061:	WC_Mult port map (I1 => X061, I2 => Coeff061, O => MultOut061, In1IW => Mult061aIW, In1FW => Mult061aFW, In2IW => Mult061bIW, In2FW => Mult061bFW);
	WC_Mult062:	WC_Mult port map (I1 => X062, I2 => Coeff062, O => MultOut062, In1IW => Mult062aIW, In1FW => Mult062aFW, In2IW => Mult062bIW, In2FW => Mult062bFW);
	WC_Mult063:	WC_Mult port map (I1 => X063, I2 => Coeff063, O => MultOut063, In1IW => Mult063aIW, In1FW => Mult063aFW, In2IW => Mult063bIW, In2FW => Mult063bFW);
	WC_Mult064:	WC_Mult port map (I1 => X064, I2 => Coeff064, O => MultOut064, In1IW => Mult064aIW, In1FW => Mult064aFW, In2IW => Mult064bIW, In2FW => Mult064bFW);
	WC_Mult065:	WC_Mult port map (I1 => X065, I2 => Coeff065, O => MultOut065, In1IW => Mult065aIW, In1FW => Mult065aFW, In2IW => Mult065bIW, In2FW => Mult065bFW);
	WC_Mult066:	WC_Mult port map (I1 => X066, I2 => Coeff066, O => MultOut066, In1IW => Mult066aIW, In1FW => Mult066aFW, In2IW => Mult066bIW, In2FW => Mult066bFW);
	WC_Mult067:	WC_Mult port map (I1 => X067, I2 => Coeff067, O => MultOut067, In1IW => Mult067aIW, In1FW => Mult067aFW, In2IW => Mult067bIW, In2FW => Mult067bFW);
	WC_Mult068:	WC_Mult port map (I1 => X068, I2 => Coeff068, O => MultOut068, In1IW => Mult068aIW, In1FW => Mult068aFW, In2IW => Mult068bIW, In2FW => Mult068bFW);
	WC_Mult069:	WC_Mult port map (I1 => X069, I2 => Coeff069, O => MultOut069, In1IW => Mult069aIW, In1FW => Mult069aFW, In2IW => Mult069bIW, In2FW => Mult069bFW);
	WC_Mult070:	WC_Mult port map (I1 => X070, I2 => Coeff070, O => MultOut070, In1IW => Mult070aIW, In1FW => Mult070aFW, In2IW => Mult070bIW, In2FW => Mult070bFW);
	WC_Mult071:	WC_Mult port map (I1 => X071, I2 => Coeff071, O => MultOut071, In1IW => Mult071aIW, In1FW => Mult071aFW, In2IW => Mult071bIW, In2FW => Mult071bFW);
	WC_Mult072:	WC_Mult port map (I1 => X072, I2 => Coeff072, O => MultOut072, In1IW => Mult072aIW, In1FW => Mult072aFW, In2IW => Mult072bIW, In2FW => Mult072bFW);
	WC_Mult073:	WC_Mult port map (I1 => X073, I2 => Coeff073, O => MultOut073, In1IW => Mult073aIW, In1FW => Mult073aFW, In2IW => Mult073bIW, In2FW => Mult073bFW);
	WC_Mult074:	WC_Mult port map (I1 => X074, I2 => Coeff074, O => MultOut074, In1IW => Mult074aIW, In1FW => Mult074aFW, In2IW => Mult074bIW, In2FW => Mult074bFW);
	WC_Mult075:	WC_Mult port map (I1 => X075, I2 => Coeff075, O => MultOut075, In1IW => Mult075aIW, In1FW => Mult075aFW, In2IW => Mult075bIW, In2FW => Mult075bFW);
	WC_Mult076:	WC_Mult port map (I1 => X076, I2 => Coeff076, O => MultOut076, In1IW => Mult076aIW, In1FW => Mult076aFW, In2IW => Mult076bIW, In2FW => Mult076bFW);
	WC_Mult077:	WC_Mult port map (I1 => X077, I2 => Coeff077, O => MultOut077, In1IW => Mult077aIW, In1FW => Mult077aFW, In2IW => Mult077bIW, In2FW => Mult077bFW);
	WC_Mult078:	WC_Mult port map (I1 => X078, I2 => Coeff078, O => MultOut078, In1IW => Mult078aIW, In1FW => Mult078aFW, In2IW => Mult078bIW, In2FW => Mult078bFW);
	WC_Mult079:	WC_Mult port map (I1 => X079, I2 => Coeff079, O => MultOut079, In1IW => Mult079aIW, In1FW => Mult079aFW, In2IW => Mult079bIW, In2FW => Mult079bFW);
	WC_Mult080:	WC_Mult port map (I1 => X080, I2 => Coeff080, O => MultOut080, In1IW => Mult080aIW, In1FW => Mult080aFW, In2IW => Mult080bIW, In2FW => Mult080bFW);
	WC_Mult081:	WC_Mult port map (I1 => X081, I2 => Coeff081, O => MultOut081, In1IW => Mult081aIW, In1FW => Mult081aFW, In2IW => Mult081bIW, In2FW => Mult081bFW);
	WC_Mult082:	WC_Mult port map (I1 => X082, I2 => Coeff082, O => MultOut082, In1IW => Mult082aIW, In1FW => Mult082aFW, In2IW => Mult082bIW, In2FW => Mult082bFW);
	WC_Mult083:	WC_Mult port map (I1 => X083, I2 => Coeff083, O => MultOut083, In1IW => Mult083aIW, In1FW => Mult083aFW, In2IW => Mult083bIW, In2FW => Mult083bFW);
	WC_Mult084:	WC_Mult port map (I1 => X084, I2 => Coeff084, O => MultOut084, In1IW => Mult084aIW, In1FW => Mult084aFW, In2IW => Mult084bIW, In2FW => Mult084bFW);
	WC_Mult085:	WC_Mult port map (I1 => X085, I2 => Coeff085, O => MultOut085, In1IW => Mult085aIW, In1FW => Mult085aFW, In2IW => Mult085bIW, In2FW => Mult085bFW);
	WC_Mult086:	WC_Mult port map (I1 => X086, I2 => Coeff086, O => MultOut086, In1IW => Mult086aIW, In1FW => Mult086aFW, In2IW => Mult086bIW, In2FW => Mult086bFW);
	WC_Mult087:	WC_Mult port map (I1 => X087, I2 => Coeff087, O => MultOut087, In1IW => Mult087aIW, In1FW => Mult087aFW, In2IW => Mult087bIW, In2FW => Mult087bFW);
	WC_Mult088:	WC_Mult port map (I1 => X088, I2 => Coeff088, O => MultOut088, In1IW => Mult088aIW, In1FW => Mult088aFW, In2IW => Mult088bIW, In2FW => Mult088bFW);
	WC_Mult089:	WC_Mult port map (I1 => X089, I2 => Coeff089, O => MultOut089, In1IW => Mult089aIW, In1FW => Mult089aFW, In2IW => Mult089bIW, In2FW => Mult089bFW);
	WC_Mult090:	WC_Mult port map (I1 => X090, I2 => Coeff090, O => MultOut090, In1IW => Mult090aIW, In1FW => Mult090aFW, In2IW => Mult090bIW, In2FW => Mult090bFW);
	WC_Mult091:	WC_Mult port map (I1 => X091, I2 => Coeff091, O => MultOut091, In1IW => Mult091aIW, In1FW => Mult091aFW, In2IW => Mult091bIW, In2FW => Mult091bFW);
	WC_Mult092:	WC_Mult port map (I1 => X092, I2 => Coeff092, O => MultOut092, In1IW => Mult092aIW, In1FW => Mult092aFW, In2IW => Mult092bIW, In2FW => Mult092bFW);
	WC_Mult093:	WC_Mult port map (I1 => X093, I2 => Coeff093, O => MultOut093, In1IW => Mult093aIW, In1FW => Mult093aFW, In2IW => Mult093bIW, In2FW => Mult093bFW);
	WC_Mult094:	WC_Mult port map (I1 => X094, I2 => Coeff094, O => MultOut094, In1IW => Mult094aIW, In1FW => Mult094aFW, In2IW => Mult094bIW, In2FW => Mult094bFW);
	WC_Mult095:	WC_Mult port map (I1 => X095, I2 => Coeff095, O => MultOut095, In1IW => Mult095aIW, In1FW => Mult095aFW, In2IW => Mult095bIW, In2FW => Mult095bFW);
	WC_Mult096:	WC_Mult port map (I1 => X096, I2 => Coeff096, O => MultOut096, In1IW => Mult096aIW, In1FW => Mult096aFW, In2IW => Mult096bIW, In2FW => Mult096bFW);
	WC_Mult097:	WC_Mult port map (I1 => X097, I2 => Coeff097, O => MultOut097, In1IW => Mult097aIW, In1FW => Mult097aFW, In2IW => Mult097bIW, In2FW => Mult097bFW);
	WC_Mult098:	WC_Mult port map (I1 => X098, I2 => Coeff098, O => MultOut098, In1IW => Mult098aIW, In1FW => Mult098aFW, In2IW => Mult098bIW, In2FW => Mult098bFW);
	WC_Mult099:	WC_Mult port map (I1 => X099, I2 => Coeff099, O => MultOut099, In1IW => Mult099aIW, In1FW => Mult099aFW, In2IW => Mult099bIW, In2FW => Mult099bFW);
	WC_Mult100:	WC_Mult port map (I1 => X100, I2 => Coeff100, O => MultOut100, In1IW => Mult100aIW, In1FW => Mult100aFW, In2IW => Mult100bIW, In2FW => Mult100bFW);
	WC_Mult101:	WC_Mult port map (I1 => X101, I2 => Coeff101, O => MultOut101, In1IW => Mult101aIW, In1FW => Mult101aFW, In2IW => Mult101bIW, In2FW => Mult101bFW);
	WC_Mult102:	WC_Mult port map (I1 => X102, I2 => Coeff102, O => MultOut102, In1IW => Mult102aIW, In1FW => Mult102aFW, In2IW => Mult102bIW, In2FW => Mult102bFW);
	WC_Mult103:	WC_Mult port map (I1 => X103, I2 => Coeff103, O => MultOut103, In1IW => Mult103aIW, In1FW => Mult103aFW, In2IW => Mult103bIW, In2FW => Mult103bFW);
	WC_Mult104:	WC_Mult port map (I1 => X104, I2 => Coeff104, O => MultOut104, In1IW => Mult104aIW, In1FW => Mult104aFW, In2IW => Mult104bIW, In2FW => Mult104bFW);
	WC_Mult105:	WC_Mult port map (I1 => X105, I2 => Coeff105, O => MultOut105, In1IW => Mult105aIW, In1FW => Mult105aFW, In2IW => Mult105bIW, In2FW => Mult105bFW);
	WC_Mult106:	WC_Mult port map (I1 => X106, I2 => Coeff106, O => MultOut106, In1IW => Mult106aIW, In1FW => Mult106aFW, In2IW => Mult106bIW, In2FW => Mult106bFW);
	WC_Mult107:	WC_Mult port map (I1 => X107, I2 => Coeff107, O => MultOut107, In1IW => Mult107aIW, In1FW => Mult107aFW, In2IW => Mult107bIW, In2FW => Mult107bFW);
	WC_Mult108:	WC_Mult port map (I1 => X108, I2 => Coeff108, O => MultOut108, In1IW => Mult108aIW, In1FW => Mult108aFW, In2IW => Mult108bIW, In2FW => Mult108bFW);
	WC_Mult109:	WC_Mult port map (I1 => X109, I2 => Coeff109, O => MultOut109, In1IW => Mult109aIW, In1FW => Mult109aFW, In2IW => Mult109bIW, In2FW => Mult109bFW);
	WC_Mult110:	WC_Mult port map (I1 => X110, I2 => Coeff110, O => MultOut110, In1IW => Mult110aIW, In1FW => Mult110aFW, In2IW => Mult110bIW, In2FW => Mult110bFW);
	WC_Mult111:	WC_Mult port map (I1 => X111, I2 => Coeff111, O => MultOut111, In1IW => Mult111aIW, In1FW => Mult111aFW, In2IW => Mult111bIW, In2FW => Mult111bFW);
	WC_Mult112:	WC_Mult port map (I1 => X112, I2 => Coeff112, O => MultOut112, In1IW => Mult112aIW, In1FW => Mult112aFW, In2IW => Mult112bIW, In2FW => Mult112bFW);
	WC_Mult113:	WC_Mult port map (I1 => X113, I2 => Coeff113, O => MultOut113, In1IW => Mult113aIW, In1FW => Mult113aFW, In2IW => Mult113bIW, In2FW => Mult113bFW);
	WC_Mult114:	WC_Mult port map (I1 => X114, I2 => Coeff114, O => MultOut114, In1IW => Mult114aIW, In1FW => Mult114aFW, In2IW => Mult114bIW, In2FW => Mult114bFW);
	WC_Mult115:	WC_Mult port map (I1 => X115, I2 => Coeff115, O => MultOut115, In1IW => Mult115aIW, In1FW => Mult115aFW, In2IW => Mult115bIW, In2FW => Mult115bFW);
	WC_Mult116:	WC_Mult port map (I1 => X116, I2 => Coeff116, O => MultOut116, In1IW => Mult116aIW, In1FW => Mult116aFW, In2IW => Mult116bIW, In2FW => Mult116bFW);
	WC_Mult117:	WC_Mult port map (I1 => X117, I2 => Coeff117, O => MultOut117, In1IW => Mult117aIW, In1FW => Mult117aFW, In2IW => Mult117bIW, In2FW => Mult117bFW);
	WC_Mult118:	WC_Mult port map (I1 => X118, I2 => Coeff118, O => MultOut118, In1IW => Mult118aIW, In1FW => Mult118aFW, In2IW => Mult118bIW, In2FW => Mult118bFW);
	WC_Mult119:	WC_Mult port map (I1 => X119, I2 => Coeff119, O => MultOut119, In1IW => Mult119aIW, In1FW => Mult119aFW, In2IW => Mult119bIW, In2FW => Mult119bFW);
	WC_Mult120:	WC_Mult port map (I1 => X120, I2 => Coeff120, O => MultOut120, In1IW => Mult120aIW, In1FW => Mult120aFW, In2IW => Mult120bIW, In2FW => Mult120bFW);
	WC_Mult121:	WC_Mult port map (I1 => X121, I2 => Coeff121, O => MultOut121, In1IW => Mult121aIW, In1FW => Mult121aFW, In2IW => Mult121bIW, In2FW => Mult121bFW);
	WC_Mult122:	WC_Mult port map (I1 => X122, I2 => Coeff122, O => MultOut122, In1IW => Mult122aIW, In1FW => Mult122aFW, In2IW => Mult122bIW, In2FW => Mult122bFW);
	WC_Mult123:	WC_Mult port map (I1 => X123, I2 => Coeff123, O => MultOut123, In1IW => Mult123aIW, In1FW => Mult123aFW, In2IW => Mult123bIW, In2FW => Mult123bFW);
	WC_Mult124:	WC_Mult port map (I1 => X124, I2 => Coeff124, O => MultOut124, In1IW => Mult124aIW, In1FW => Mult124aFW, In2IW => Mult124bIW, In2FW => Mult124bFW);
	WC_Mult125:	WC_Mult port map (I1 => X125, I2 => Coeff125, O => MultOut125, In1IW => Mult125aIW, In1FW => Mult125aFW, In2IW => Mult125bIW, In2FW => Mult125bFW);
	WC_Mult126:	WC_Mult port map (I1 => X126, I2 => Coeff126, O => MultOut126, In1IW => Mult126aIW, In1FW => Mult126aFW, In2IW => Mult126bIW, In2FW => Mult126bFW);
	WC_Mult127:	WC_Mult port map (I1 => X127, I2 => Coeff127, O => MultOut127, In1IW => Mult127aIW, In1FW => Mult127aFW, In2IW => Mult127bIW, In2FW => Mult127bFW);
	WC_Mult128:	WC_Mult port map (I1 => X128, I2 => Coeff128, O => MultOut128, In1IW => Mult128aIW, In1FW => Mult128aFW, In2IW => Mult128bIW, In2FW => Mult128bFW);
	WC_Mult129:	WC_Mult port map (I1 => X129, I2 => Coeff129, O => MultOut129, In1IW => Mult129aIW, In1FW => Mult129aFW, In2IW => Mult129bIW, In2FW => Mult129bFW);
	WC_Mult130:	WC_Mult port map (I1 => X130, I2 => Coeff130, O => MultOut130, In1IW => Mult130aIW, In1FW => Mult130aFW, In2IW => Mult130bIW, In2FW => Mult130bFW);
	WC_Mult131:	WC_Mult port map (I1 => X131, I2 => Coeff131, O => MultOut131, In1IW => Mult131aIW, In1FW => Mult131aFW, In2IW => Mult131bIW, In2FW => Mult131bFW);
	WC_Mult132:	WC_Mult port map (I1 => X132, I2 => Coeff132, O => MultOut132, In1IW => Mult132aIW, In1FW => Mult132aFW, In2IW => Mult132bIW, In2FW => Mult132bFW);
	WC_Mult133:	WC_Mult port map (I1 => X133, I2 => Coeff133, O => MultOut133, In1IW => Mult133aIW, In1FW => Mult133aFW, In2IW => Mult133bIW, In2FW => Mult133bFW);
	WC_Mult134:	WC_Mult port map (I1 => X134, I2 => Coeff134, O => MultOut134, In1IW => Mult134aIW, In1FW => Mult134aFW, In2IW => Mult134bIW, In2FW => Mult134bFW);
	WC_Mult135:	WC_Mult port map (I1 => X135, I2 => Coeff135, O => MultOut135, In1IW => Mult135aIW, In1FW => Mult135aFW, In2IW => Mult135bIW, In2FW => Mult135bFW);
	WC_Mult136:	WC_Mult port map (I1 => X136, I2 => Coeff136, O => MultOut136, In1IW => Mult136aIW, In1FW => Mult136aFW, In2IW => Mult136bIW, In2FW => Mult136bFW);
	WC_Mult137:	WC_Mult port map (I1 => X137, I2 => Coeff137, O => MultOut137, In1IW => Mult137aIW, In1FW => Mult137aFW, In2IW => Mult137bIW, In2FW => Mult137bFW);
	WC_Mult138:	WC_Mult port map (I1 => X138, I2 => Coeff138, O => MultOut138, In1IW => Mult138aIW, In1FW => Mult138aFW, In2IW => Mult138bIW, In2FW => Mult138bFW);
	WC_Mult139:	WC_Mult port map (I1 => X139, I2 => Coeff139, O => MultOut139, In1IW => Mult139aIW, In1FW => Mult139aFW, In2IW => Mult139bIW, In2FW => Mult139bFW);
	WC_Mult140:	WC_Mult port map (I1 => X140, I2 => Coeff140, O => MultOut140, In1IW => Mult140aIW, In1FW => Mult140aFW, In2IW => Mult140bIW, In2FW => Mult140bFW);
	WC_Mult141:	WC_Mult port map (I1 => X141, I2 => Coeff141, O => MultOut141, In1IW => Mult141aIW, In1FW => Mult141aFW, In2IW => Mult141bIW, In2FW => Mult141bFW);
	WC_Mult142:	WC_Mult port map (I1 => X142, I2 => Coeff142, O => MultOut142, In1IW => Mult142aIW, In1FW => Mult142aFW, In2IW => Mult142bIW, In2FW => Mult142bFW);
	WC_Mult143:	WC_Mult port map (I1 => X143, I2 => Coeff143, O => MultOut143, In1IW => Mult143aIW, In1FW => Mult143aFW, In2IW => Mult143bIW, In2FW => Mult143bFW);
	WC_Mult144:	WC_Mult port map (I1 => X144, I2 => Coeff144, O => MultOut144, In1IW => Mult144aIW, In1FW => Mult144aFW, In2IW => Mult144bIW, In2FW => Mult144bFW);
	WC_Mult145:	WC_Mult port map (I1 => X145, I2 => Coeff145, O => MultOut145, In1IW => Mult145aIW, In1FW => Mult145aFW, In2IW => Mult145bIW, In2FW => Mult145bFW);
	WC_Mult146:	WC_Mult port map (I1 => X146, I2 => Coeff146, O => MultOut146, In1IW => Mult146aIW, In1FW => Mult146aFW, In2IW => Mult146bIW, In2FW => Mult146bFW);
	WC_Mult147:	WC_Mult port map (I1 => X147, I2 => Coeff147, O => MultOut147, In1IW => Mult147aIW, In1FW => Mult147aFW, In2IW => Mult147bIW, In2FW => Mult147bFW);
	WC_Mult148:	WC_Mult port map (I1 => X148, I2 => Coeff148, O => MultOut148, In1IW => Mult148aIW, In1FW => Mult148aFW, In2IW => Mult148bIW, In2FW => Mult148bFW);
	WC_Mult149:	WC_Mult port map (I1 => X149, I2 => Coeff149, O => MultOut149, In1IW => Mult149aIW, In1FW => Mult149aFW, In2IW => Mult149bIW, In2FW => Mult149bFW);
	WC_Mult150:	WC_Mult port map (I1 => X150, I2 => Coeff150, O => MultOut150, In1IW => Mult150aIW, In1FW => Mult150aFW, In2IW => Mult150bIW, In2FW => Mult150bFW);

	
	-- Adders
	WC_Adder000:	WC_AddSub port map (I1 => Y000, I2 => MultOut000, O => Y001, In1IW => Add000aIW, In1FW => Add000aFW, In2IW => Add000bIW, In2FW => Add000bFW);
	WC_Adder001:	WC_AddSub port map (I1 => Y001, I2 => MultOut001, O => Y002, In1IW => Add001aIW, In1FW => Add001aFW, In2IW => Add001bIW, In2FW => Add001bFW);
	WC_Adder002:	WC_AddSub port map (I1 => Y002, I2 => MultOut002, O => Y003, In1IW => Add002aIW, In1FW => Add002aFW, In2IW => Add002bIW, In2FW => Add002bFW);
	WC_Adder003:	WC_AddSub port map (I1 => Y003, I2 => MultOut003, O => Y004, In1IW => Add003aIW, In1FW => Add003aFW, In2IW => Add003bIW, In2FW => Add003bFW);
	WC_Adder004:	WC_AddSub port map (I1 => Y004, I2 => MultOut004, O => Y005, In1IW => Add004aIW, In1FW => Add004aFW, In2IW => Add004bIW, In2FW => Add004bFW);
	WC_Adder005:	WC_AddSub port map (I1 => Y005, I2 => MultOut005, O => Y006, In1IW => Add005aIW, In1FW => Add005aFW, In2IW => Add005bIW, In2FW => Add005bFW);
	WC_Adder006:	WC_AddSub port map (I1 => Y006, I2 => MultOut006, O => Y007, In1IW => Add006aIW, In1FW => Add006aFW, In2IW => Add006bIW, In2FW => Add006bFW);
	WC_Adder007:	WC_AddSub port map (I1 => Y007, I2 => MultOut007, O => Y008, In1IW => Add007aIW, In1FW => Add007aFW, In2IW => Add007bIW, In2FW => Add007bFW);
	WC_Adder008:	WC_AddSub port map (I1 => Y008, I2 => MultOut008, O => Y009, In1IW => Add008aIW, In1FW => Add008aFW, In2IW => Add008bIW, In2FW => Add008bFW);
	WC_Adder009:	WC_AddSub port map (I1 => Y009, I2 => MultOut009, O => Y010, In1IW => Add009aIW, In1FW => Add009aFW, In2IW => Add009bIW, In2FW => Add009bFW);
	WC_Adder010:	WC_AddSub port map (I1 => Y010, I2 => MultOut010, O => Y011, In1IW => Add010aIW, In1FW => Add010aFW, In2IW => Add010bIW, In2FW => Add010bFW);
	WC_Adder011:	WC_AddSub port map (I1 => Y011, I2 => MultOut011, O => Y012, In1IW => Add011aIW, In1FW => Add011aFW, In2IW => Add011bIW, In2FW => Add011bFW);
	WC_Adder012:	WC_AddSub port map (I1 => Y012, I2 => MultOut012, O => Y013, In1IW => Add012aIW, In1FW => Add012aFW, In2IW => Add012bIW, In2FW => Add012bFW);
	WC_Adder013:	WC_AddSub port map (I1 => Y013, I2 => MultOut013, O => Y014, In1IW => Add013aIW, In1FW => Add013aFW, In2IW => Add013bIW, In2FW => Add013bFW);
	WC_Adder014:	WC_AddSub port map (I1 => Y014, I2 => MultOut014, O => Y015, In1IW => Add014aIW, In1FW => Add014aFW, In2IW => Add014bIW, In2FW => Add014bFW);
	WC_Adder015:	WC_AddSub port map (I1 => Y015, I2 => MultOut015, O => Y016, In1IW => Add015aIW, In1FW => Add015aFW, In2IW => Add015bIW, In2FW => Add015bFW);
	WC_Adder016:	WC_AddSub port map (I1 => Y016, I2 => MultOut016, O => Y017, In1IW => Add016aIW, In1FW => Add016aFW, In2IW => Add016bIW, In2FW => Add016bFW);
	WC_Adder017:	WC_AddSub port map (I1 => Y017, I2 => MultOut017, O => Y018, In1IW => Add017aIW, In1FW => Add017aFW, In2IW => Add017bIW, In2FW => Add017bFW);
	WC_Adder018:	WC_AddSub port map (I1 => Y018, I2 => MultOut018, O => Y019, In1IW => Add018aIW, In1FW => Add018aFW, In2IW => Add018bIW, In2FW => Add018bFW);
	WC_Adder019:	WC_AddSub port map (I1 => Y019, I2 => MultOut019, O => Y020, In1IW => Add019aIW, In1FW => Add019aFW, In2IW => Add019bIW, In2FW => Add019bFW);
	WC_Adder020:	WC_AddSub port map (I1 => Y020, I2 => MultOut020, O => Y021, In1IW => Add020aIW, In1FW => Add020aFW, In2IW => Add020bIW, In2FW => Add020bFW);
	WC_Adder021:	WC_AddSub port map (I1 => Y021, I2 => MultOut021, O => Y022, In1IW => Add021aIW, In1FW => Add021aFW, In2IW => Add021bIW, In2FW => Add021bFW);
	WC_Adder022:	WC_AddSub port map (I1 => Y022, I2 => MultOut022, O => Y023, In1IW => Add022aIW, In1FW => Add022aFW, In2IW => Add022bIW, In2FW => Add022bFW);
	WC_Adder023:	WC_AddSub port map (I1 => Y023, I2 => MultOut023, O => Y024, In1IW => Add023aIW, In1FW => Add023aFW, In2IW => Add023bIW, In2FW => Add023bFW);
	WC_Adder024:	WC_AddSub port map (I1 => Y024, I2 => MultOut024, O => Y025, In1IW => Add024aIW, In1FW => Add024aFW, In2IW => Add024bIW, In2FW => Add024bFW);
	WC_Adder025:	WC_AddSub port map (I1 => Y025, I2 => MultOut025, O => Y026, In1IW => Add025aIW, In1FW => Add025aFW, In2IW => Add025bIW, In2FW => Add025bFW);
	WC_Adder026:	WC_AddSub port map (I1 => Y026, I2 => MultOut026, O => Y027, In1IW => Add026aIW, In1FW => Add026aFW, In2IW => Add026bIW, In2FW => Add026bFW);
	WC_Adder027:	WC_AddSub port map (I1 => Y027, I2 => MultOut027, O => Y028, In1IW => Add027aIW, In1FW => Add027aFW, In2IW => Add027bIW, In2FW => Add027bFW);
	WC_Adder028:	WC_AddSub port map (I1 => Y028, I2 => MultOut028, O => Y029, In1IW => Add028aIW, In1FW => Add028aFW, In2IW => Add028bIW, In2FW => Add028bFW);
	WC_Adder029:	WC_AddSub port map (I1 => Y029, I2 => MultOut029, O => Y030, In1IW => Add029aIW, In1FW => Add029aFW, In2IW => Add029bIW, In2FW => Add029bFW);
	WC_Adder030:	WC_AddSub port map (I1 => Y030, I2 => MultOut030, O => Y031, In1IW => Add030aIW, In1FW => Add030aFW, In2IW => Add030bIW, In2FW => Add030bFW);
	WC_Adder031:	WC_AddSub port map (I1 => Y031, I2 => MultOut031, O => Y032, In1IW => Add031aIW, In1FW => Add031aFW, In2IW => Add031bIW, In2FW => Add031bFW);
	WC_Adder032:	WC_AddSub port map (I1 => Y032, I2 => MultOut032, O => Y033, In1IW => Add032aIW, In1FW => Add032aFW, In2IW => Add032bIW, In2FW => Add032bFW);
	WC_Adder033:	WC_AddSub port map (I1 => Y033, I2 => MultOut033, O => Y034, In1IW => Add033aIW, In1FW => Add033aFW, In2IW => Add033bIW, In2FW => Add033bFW);
	WC_Adder034:	WC_AddSub port map (I1 => Y034, I2 => MultOut034, O => Y035, In1IW => Add034aIW, In1FW => Add034aFW, In2IW => Add034bIW, In2FW => Add034bFW);
	WC_Adder035:	WC_AddSub port map (I1 => Y035, I2 => MultOut035, O => Y036, In1IW => Add035aIW, In1FW => Add035aFW, In2IW => Add035bIW, In2FW => Add035bFW);
	WC_Adder036:	WC_AddSub port map (I1 => Y036, I2 => MultOut036, O => Y037, In1IW => Add036aIW, In1FW => Add036aFW, In2IW => Add036bIW, In2FW => Add036bFW);
	WC_Adder037:	WC_AddSub port map (I1 => Y037, I2 => MultOut037, O => Y038, In1IW => Add037aIW, In1FW => Add037aFW, In2IW => Add037bIW, In2FW => Add037bFW);
	WC_Adder038:	WC_AddSub port map (I1 => Y038, I2 => MultOut038, O => Y039, In1IW => Add038aIW, In1FW => Add038aFW, In2IW => Add038bIW, In2FW => Add038bFW);
	WC_Adder039:	WC_AddSub port map (I1 => Y039, I2 => MultOut039, O => Y040, In1IW => Add039aIW, In1FW => Add039aFW, In2IW => Add039bIW, In2FW => Add039bFW);
	WC_Adder040:	WC_AddSub port map (I1 => Y040, I2 => MultOut040, O => Y041, In1IW => Add040aIW, In1FW => Add040aFW, In2IW => Add040bIW, In2FW => Add040bFW);
	WC_Adder041:	WC_AddSub port map (I1 => Y041, I2 => MultOut041, O => Y042, In1IW => Add041aIW, In1FW => Add041aFW, In2IW => Add041bIW, In2FW => Add041bFW);
	WC_Adder042:	WC_AddSub port map (I1 => Y042, I2 => MultOut042, O => Y043, In1IW => Add042aIW, In1FW => Add042aFW, In2IW => Add042bIW, In2FW => Add042bFW);
	WC_Adder043:	WC_AddSub port map (I1 => Y043, I2 => MultOut043, O => Y044, In1IW => Add043aIW, In1FW => Add043aFW, In2IW => Add043bIW, In2FW => Add043bFW);
	WC_Adder044:	WC_AddSub port map (I1 => Y044, I2 => MultOut044, O => Y045, In1IW => Add044aIW, In1FW => Add044aFW, In2IW => Add044bIW, In2FW => Add044bFW);
	WC_Adder045:	WC_AddSub port map (I1 => Y045, I2 => MultOut045, O => Y046, In1IW => Add045aIW, In1FW => Add045aFW, In2IW => Add045bIW, In2FW => Add045bFW);
	WC_Adder046:	WC_AddSub port map (I1 => Y046, I2 => MultOut046, O => Y047, In1IW => Add046aIW, In1FW => Add046aFW, In2IW => Add046bIW, In2FW => Add046bFW);
	WC_Adder047:	WC_AddSub port map (I1 => Y047, I2 => MultOut047, O => Y048, In1IW => Add047aIW, In1FW => Add047aFW, In2IW => Add047bIW, In2FW => Add047bFW);
	WC_Adder048:	WC_AddSub port map (I1 => Y048, I2 => MultOut048, O => Y049, In1IW => Add048aIW, In1FW => Add048aFW, In2IW => Add048bIW, In2FW => Add048bFW);
	WC_Adder049:	WC_AddSub port map (I1 => Y049, I2 => MultOut049, O => Y050, In1IW => Add049aIW, In1FW => Add049aFW, In2IW => Add049bIW, In2FW => Add049bFW);
	WC_Adder050:	WC_AddSub port map (I1 => Y050, I2 => MultOut050, O => Y051, In1IW => Add050aIW, In1FW => Add050aFW, In2IW => Add050bIW, In2FW => Add050bFW);
	WC_Adder051:	WC_AddSub port map (I1 => Y051, I2 => MultOut051, O => Y052, In1IW => Add051aIW, In1FW => Add051aFW, In2IW => Add051bIW, In2FW => Add051bFW);
	WC_Adder052:	WC_AddSub port map (I1 => Y052, I2 => MultOut052, O => Y053, In1IW => Add052aIW, In1FW => Add052aFW, In2IW => Add052bIW, In2FW => Add052bFW);
	WC_Adder053:	WC_AddSub port map (I1 => Y053, I2 => MultOut053, O => Y054, In1IW => Add053aIW, In1FW => Add053aFW, In2IW => Add053bIW, In2FW => Add053bFW);
	WC_Adder054:	WC_AddSub port map (I1 => Y054, I2 => MultOut054, O => Y055, In1IW => Add054aIW, In1FW => Add054aFW, In2IW => Add054bIW, In2FW => Add054bFW);
	WC_Adder055:	WC_AddSub port map (I1 => Y055, I2 => MultOut055, O => Y056, In1IW => Add055aIW, In1FW => Add055aFW, In2IW => Add055bIW, In2FW => Add055bFW);
	WC_Adder056:	WC_AddSub port map (I1 => Y056, I2 => MultOut056, O => Y057, In1IW => Add056aIW, In1FW => Add056aFW, In2IW => Add056bIW, In2FW => Add056bFW);
	WC_Adder057:	WC_AddSub port map (I1 => Y057, I2 => MultOut057, O => Y058, In1IW => Add057aIW, In1FW => Add057aFW, In2IW => Add057bIW, In2FW => Add057bFW);
	WC_Adder058:	WC_AddSub port map (I1 => Y058, I2 => MultOut058, O => Y059, In1IW => Add058aIW, In1FW => Add058aFW, In2IW => Add058bIW, In2FW => Add058bFW);
	WC_Adder059:	WC_AddSub port map (I1 => Y059, I2 => MultOut059, O => Y060, In1IW => Add059aIW, In1FW => Add059aFW, In2IW => Add059bIW, In2FW => Add059bFW);
	WC_Adder060:	WC_AddSub port map (I1 => Y060, I2 => MultOut060, O => Y061, In1IW => Add060aIW, In1FW => Add060aFW, In2IW => Add060bIW, In2FW => Add060bFW);
	WC_Adder061:	WC_AddSub port map (I1 => Y061, I2 => MultOut061, O => Y062, In1IW => Add061aIW, In1FW => Add061aFW, In2IW => Add061bIW, In2FW => Add061bFW);
	WC_Adder062:	WC_AddSub port map (I1 => Y062, I2 => MultOut062, O => Y063, In1IW => Add062aIW, In1FW => Add062aFW, In2IW => Add062bIW, In2FW => Add062bFW);
	WC_Adder063:	WC_AddSub port map (I1 => Y063, I2 => MultOut063, O => Y064, In1IW => Add063aIW, In1FW => Add063aFW, In2IW => Add063bIW, In2FW => Add063bFW);
	WC_Adder064:	WC_AddSub port map (I1 => Y064, I2 => MultOut064, O => Y065, In1IW => Add064aIW, In1FW => Add064aFW, In2IW => Add064bIW, In2FW => Add064bFW);
	WC_Adder065:	WC_AddSub port map (I1 => Y065, I2 => MultOut065, O => Y066, In1IW => Add065aIW, In1FW => Add065aFW, In2IW => Add065bIW, In2FW => Add065bFW);
	WC_Adder066:	WC_AddSub port map (I1 => Y066, I2 => MultOut066, O => Y067, In1IW => Add066aIW, In1FW => Add066aFW, In2IW => Add066bIW, In2FW => Add066bFW);
	WC_Adder067:	WC_AddSub port map (I1 => Y067, I2 => MultOut067, O => Y068, In1IW => Add067aIW, In1FW => Add067aFW, In2IW => Add067bIW, In2FW => Add067bFW);
	WC_Adder068:	WC_AddSub port map (I1 => Y068, I2 => MultOut068, O => Y069, In1IW => Add068aIW, In1FW => Add068aFW, In2IW => Add068bIW, In2FW => Add068bFW);
	WC_Adder069:	WC_AddSub port map (I1 => Y069, I2 => MultOut069, O => Y070, In1IW => Add069aIW, In1FW => Add069aFW, In2IW => Add069bIW, In2FW => Add069bFW);
	WC_Adder070:	WC_AddSub port map (I1 => Y070, I2 => MultOut070, O => Y071, In1IW => Add070aIW, In1FW => Add070aFW, In2IW => Add070bIW, In2FW => Add070bFW);
	WC_Adder071:	WC_AddSub port map (I1 => Y071, I2 => MultOut071, O => Y072, In1IW => Add071aIW, In1FW => Add071aFW, In2IW => Add071bIW, In2FW => Add071bFW);
	WC_Adder072:	WC_AddSub port map (I1 => Y072, I2 => MultOut072, O => Y073, In1IW => Add072aIW, In1FW => Add072aFW, In2IW => Add072bIW, In2FW => Add072bFW);
	WC_Adder073:	WC_AddSub port map (I1 => Y073, I2 => MultOut073, O => Y074, In1IW => Add073aIW, In1FW => Add073aFW, In2IW => Add073bIW, In2FW => Add073bFW);
	WC_Adder074:	WC_AddSub port map (I1 => Y074, I2 => MultOut074, O => Y075, In1IW => Add074aIW, In1FW => Add074aFW, In2IW => Add074bIW, In2FW => Add074bFW);
	WC_Adder075:	WC_AddSub port map (I1 => Y075, I2 => MultOut075, O => Y076, In1IW => Add075aIW, In1FW => Add075aFW, In2IW => Add075bIW, In2FW => Add075bFW);
	WC_Adder076:	WC_AddSub port map (I1 => Y076, I2 => MultOut076, O => Y077, In1IW => Add076aIW, In1FW => Add076aFW, In2IW => Add076bIW, In2FW => Add076bFW);
	WC_Adder077:	WC_AddSub port map (I1 => Y077, I2 => MultOut077, O => Y078, In1IW => Add077aIW, In1FW => Add077aFW, In2IW => Add077bIW, In2FW => Add077bFW);
	WC_Adder078:	WC_AddSub port map (I1 => Y078, I2 => MultOut078, O => Y079, In1IW => Add078aIW, In1FW => Add078aFW, In2IW => Add078bIW, In2FW => Add078bFW);
	WC_Adder079:	WC_AddSub port map (I1 => Y079, I2 => MultOut079, O => Y080, In1IW => Add079aIW, In1FW => Add079aFW, In2IW => Add079bIW, In2FW => Add079bFW);
	WC_Adder080:	WC_AddSub port map (I1 => Y080, I2 => MultOut080, O => Y081, In1IW => Add080aIW, In1FW => Add080aFW, In2IW => Add080bIW, In2FW => Add080bFW);
	WC_Adder081:	WC_AddSub port map (I1 => Y081, I2 => MultOut081, O => Y082, In1IW => Add081aIW, In1FW => Add081aFW, In2IW => Add081bIW, In2FW => Add081bFW);
	WC_Adder082:	WC_AddSub port map (I1 => Y082, I2 => MultOut082, O => Y083, In1IW => Add082aIW, In1FW => Add082aFW, In2IW => Add082bIW, In2FW => Add082bFW);
	WC_Adder083:	WC_AddSub port map (I1 => Y083, I2 => MultOut083, O => Y084, In1IW => Add083aIW, In1FW => Add083aFW, In2IW => Add083bIW, In2FW => Add083bFW);
	WC_Adder084:	WC_AddSub port map (I1 => Y084, I2 => MultOut084, O => Y085, In1IW => Add084aIW, In1FW => Add084aFW, In2IW => Add084bIW, In2FW => Add084bFW);
	WC_Adder085:	WC_AddSub port map (I1 => Y085, I2 => MultOut085, O => Y086, In1IW => Add085aIW, In1FW => Add085aFW, In2IW => Add085bIW, In2FW => Add085bFW);
	WC_Adder086:	WC_AddSub port map (I1 => Y086, I2 => MultOut086, O => Y087, In1IW => Add086aIW, In1FW => Add086aFW, In2IW => Add086bIW, In2FW => Add086bFW);
	WC_Adder087:	WC_AddSub port map (I1 => Y087, I2 => MultOut087, O => Y088, In1IW => Add087aIW, In1FW => Add087aFW, In2IW => Add087bIW, In2FW => Add087bFW);
	WC_Adder088:	WC_AddSub port map (I1 => Y088, I2 => MultOut088, O => Y089, In1IW => Add088aIW, In1FW => Add088aFW, In2IW => Add088bIW, In2FW => Add088bFW);
	WC_Adder089:	WC_AddSub port map (I1 => Y089, I2 => MultOut089, O => Y090, In1IW => Add089aIW, In1FW => Add089aFW, In2IW => Add089bIW, In2FW => Add089bFW);
	WC_Adder090:	WC_AddSub port map (I1 => Y090, I2 => MultOut090, O => Y091, In1IW => Add090aIW, In1FW => Add090aFW, In2IW => Add090bIW, In2FW => Add090bFW);
	WC_Adder091:	WC_AddSub port map (I1 => Y091, I2 => MultOut091, O => Y092, In1IW => Add091aIW, In1FW => Add091aFW, In2IW => Add091bIW, In2FW => Add091bFW);
	WC_Adder092:	WC_AddSub port map (I1 => Y092, I2 => MultOut092, O => Y093, In1IW => Add092aIW, In1FW => Add092aFW, In2IW => Add092bIW, In2FW => Add092bFW);
	WC_Adder093:	WC_AddSub port map (I1 => Y093, I2 => MultOut093, O => Y094, In1IW => Add093aIW, In1FW => Add093aFW, In2IW => Add093bIW, In2FW => Add093bFW);
	WC_Adder094:	WC_AddSub port map (I1 => Y094, I2 => MultOut094, O => Y095, In1IW => Add094aIW, In1FW => Add094aFW, In2IW => Add094bIW, In2FW => Add094bFW);
	WC_Adder095:	WC_AddSub port map (I1 => Y095, I2 => MultOut095, O => Y096, In1IW => Add095aIW, In1FW => Add095aFW, In2IW => Add095bIW, In2FW => Add095bFW);
	WC_Adder096:	WC_AddSub port map (I1 => Y096, I2 => MultOut096, O => Y097, In1IW => Add096aIW, In1FW => Add096aFW, In2IW => Add096bIW, In2FW => Add096bFW);
	WC_Adder097:	WC_AddSub port map (I1 => Y097, I2 => MultOut097, O => Y098, In1IW => Add097aIW, In1FW => Add097aFW, In2IW => Add097bIW, In2FW => Add097bFW);
	WC_Adder098:	WC_AddSub port map (I1 => Y098, I2 => MultOut098, O => Y099, In1IW => Add098aIW, In1FW => Add098aFW, In2IW => Add098bIW, In2FW => Add098bFW);
	WC_Adder099:	WC_AddSub port map (I1 => Y099, I2 => MultOut099, O => Y100, In1IW => Add099aIW, In1FW => Add099aFW, In2IW => Add099bIW, In2FW => Add099bFW);
	WC_Adder100:	WC_AddSub port map (I1 => Y100, I2 => MultOut100, O => Y101, In1IW => Add100aIW, In1FW => Add100aFW, In2IW => Add100bIW, In2FW => Add100bFW);
	WC_Adder101:	WC_AddSub port map (I1 => Y101, I2 => MultOut101, O => Y102, In1IW => Add101aIW, In1FW => Add101aFW, In2IW => Add101bIW, In2FW => Add101bFW);
	WC_Adder102:	WC_AddSub port map (I1 => Y102, I2 => MultOut102, O => Y103, In1IW => Add102aIW, In1FW => Add102aFW, In2IW => Add102bIW, In2FW => Add102bFW);
	WC_Adder103:	WC_AddSub port map (I1 => Y103, I2 => MultOut103, O => Y104, In1IW => Add103aIW, In1FW => Add103aFW, In2IW => Add103bIW, In2FW => Add103bFW);
	WC_Adder104:	WC_AddSub port map (I1 => Y104, I2 => MultOut104, O => Y105, In1IW => Add104aIW, In1FW => Add104aFW, In2IW => Add104bIW, In2FW => Add104bFW);
	WC_Adder105:	WC_AddSub port map (I1 => Y105, I2 => MultOut105, O => Y106, In1IW => Add105aIW, In1FW => Add105aFW, In2IW => Add105bIW, In2FW => Add105bFW);
	WC_Adder106:	WC_AddSub port map (I1 => Y106, I2 => MultOut106, O => Y107, In1IW => Add106aIW, In1FW => Add106aFW, In2IW => Add106bIW, In2FW => Add106bFW);
	WC_Adder107:	WC_AddSub port map (I1 => Y107, I2 => MultOut107, O => Y108, In1IW => Add107aIW, In1FW => Add107aFW, In2IW => Add107bIW, In2FW => Add107bFW);
	WC_Adder108:	WC_AddSub port map (I1 => Y108, I2 => MultOut108, O => Y109, In1IW => Add108aIW, In1FW => Add108aFW, In2IW => Add108bIW, In2FW => Add108bFW);
	WC_Adder109:	WC_AddSub port map (I1 => Y109, I2 => MultOut109, O => Y110, In1IW => Add109aIW, In1FW => Add109aFW, In2IW => Add109bIW, In2FW => Add109bFW);
	WC_Adder110:	WC_AddSub port map (I1 => Y110, I2 => MultOut110, O => Y111, In1IW => Add110aIW, In1FW => Add110aFW, In2IW => Add110bIW, In2FW => Add110bFW);
	WC_Adder111:	WC_AddSub port map (I1 => Y111, I2 => MultOut111, O => Y112, In1IW => Add111aIW, In1FW => Add111aFW, In2IW => Add111bIW, In2FW => Add111bFW);
	WC_Adder112:	WC_AddSub port map (I1 => Y112, I2 => MultOut112, O => Y113, In1IW => Add112aIW, In1FW => Add112aFW, In2IW => Add112bIW, In2FW => Add112bFW);
	WC_Adder113:	WC_AddSub port map (I1 => Y113, I2 => MultOut113, O => Y114, In1IW => Add113aIW, In1FW => Add113aFW, In2IW => Add113bIW, In2FW => Add113bFW);
	WC_Adder114:	WC_AddSub port map (I1 => Y114, I2 => MultOut114, O => Y115, In1IW => Add114aIW, In1FW => Add114aFW, In2IW => Add114bIW, In2FW => Add114bFW);
	WC_Adder115:	WC_AddSub port map (I1 => Y115, I2 => MultOut115, O => Y116, In1IW => Add115aIW, In1FW => Add115aFW, In2IW => Add115bIW, In2FW => Add115bFW);
	WC_Adder116:	WC_AddSub port map (I1 => Y116, I2 => MultOut116, O => Y117, In1IW => Add116aIW, In1FW => Add116aFW, In2IW => Add116bIW, In2FW => Add116bFW);
	WC_Adder117:	WC_AddSub port map (I1 => Y117, I2 => MultOut117, O => Y118, In1IW => Add117aIW, In1FW => Add117aFW, In2IW => Add117bIW, In2FW => Add117bFW);
	WC_Adder118:	WC_AddSub port map (I1 => Y118, I2 => MultOut118, O => Y119, In1IW => Add118aIW, In1FW => Add118aFW, In2IW => Add118bIW, In2FW => Add118bFW);
	WC_Adder119:	WC_AddSub port map (I1 => Y119, I2 => MultOut119, O => Y120, In1IW => Add119aIW, In1FW => Add119aFW, In2IW => Add119bIW, In2FW => Add119bFW);
	WC_Adder120:	WC_AddSub port map (I1 => Y120, I2 => MultOut120, O => Y121, In1IW => Add120aIW, In1FW => Add120aFW, In2IW => Add120bIW, In2FW => Add120bFW);
	WC_Adder121:	WC_AddSub port map (I1 => Y121, I2 => MultOut121, O => Y122, In1IW => Add121aIW, In1FW => Add121aFW, In2IW => Add121bIW, In2FW => Add121bFW);
	WC_Adder122:	WC_AddSub port map (I1 => Y122, I2 => MultOut122, O => Y123, In1IW => Add122aIW, In1FW => Add122aFW, In2IW => Add122bIW, In2FW => Add122bFW);
	WC_Adder123:	WC_AddSub port map (I1 => Y123, I2 => MultOut123, O => Y124, In1IW => Add123aIW, In1FW => Add123aFW, In2IW => Add123bIW, In2FW => Add123bFW);
	WC_Adder124:	WC_AddSub port map (I1 => Y124, I2 => MultOut124, O => Y125, In1IW => Add124aIW, In1FW => Add124aFW, In2IW => Add124bIW, In2FW => Add124bFW);
	WC_Adder125:	WC_AddSub port map (I1 => Y125, I2 => MultOut125, O => Y126, In1IW => Add125aIW, In1FW => Add125aFW, In2IW => Add125bIW, In2FW => Add125bFW);
	WC_Adder126:	WC_AddSub port map (I1 => Y126, I2 => MultOut126, O => Y127, In1IW => Add126aIW, In1FW => Add126aFW, In2IW => Add126bIW, In2FW => Add126bFW);
	WC_Adder127:	WC_AddSub port map (I1 => Y127, I2 => MultOut127, O => Y128, In1IW => Add127aIW, In1FW => Add127aFW, In2IW => Add127bIW, In2FW => Add127bFW);
	WC_Adder128:	WC_AddSub port map (I1 => Y128, I2 => MultOut128, O => Y129, In1IW => Add128aIW, In1FW => Add128aFW, In2IW => Add128bIW, In2FW => Add128bFW);
	WC_Adder129:	WC_AddSub port map (I1 => Y129, I2 => MultOut129, O => Y130, In1IW => Add129aIW, In1FW => Add129aFW, In2IW => Add129bIW, In2FW => Add129bFW);
	WC_Adder130:	WC_AddSub port map (I1 => Y130, I2 => MultOut130, O => Y131, In1IW => Add130aIW, In1FW => Add130aFW, In2IW => Add130bIW, In2FW => Add130bFW);
	WC_Adder131:	WC_AddSub port map (I1 => Y131, I2 => MultOut131, O => Y132, In1IW => Add131aIW, In1FW => Add131aFW, In2IW => Add131bIW, In2FW => Add131bFW);
	WC_Adder132:	WC_AddSub port map (I1 => Y132, I2 => MultOut132, O => Y133, In1IW => Add132aIW, In1FW => Add132aFW, In2IW => Add132bIW, In2FW => Add132bFW);
	WC_Adder133:	WC_AddSub port map (I1 => Y133, I2 => MultOut133, O => Y134, In1IW => Add133aIW, In1FW => Add133aFW, In2IW => Add133bIW, In2FW => Add133bFW);
	WC_Adder134:	WC_AddSub port map (I1 => Y134, I2 => MultOut134, O => Y135, In1IW => Add134aIW, In1FW => Add134aFW, In2IW => Add134bIW, In2FW => Add134bFW);
	WC_Adder135:	WC_AddSub port map (I1 => Y135, I2 => MultOut135, O => Y136, In1IW => Add135aIW, In1FW => Add135aFW, In2IW => Add135bIW, In2FW => Add135bFW);
	WC_Adder136:	WC_AddSub port map (I1 => Y136, I2 => MultOut136, O => Y137, In1IW => Add136aIW, In1FW => Add136aFW, In2IW => Add136bIW, In2FW => Add136bFW);
	WC_Adder137:	WC_AddSub port map (I1 => Y137, I2 => MultOut137, O => Y138, In1IW => Add137aIW, In1FW => Add137aFW, In2IW => Add137bIW, In2FW => Add137bFW);
	WC_Adder138:	WC_AddSub port map (I1 => Y138, I2 => MultOut138, O => Y139, In1IW => Add138aIW, In1FW => Add138aFW, In2IW => Add138bIW, In2FW => Add138bFW);
	WC_Adder139:	WC_AddSub port map (I1 => Y139, I2 => MultOut139, O => Y140, In1IW => Add139aIW, In1FW => Add139aFW, In2IW => Add139bIW, In2FW => Add139bFW);
	WC_Adder140:	WC_AddSub port map (I1 => Y140, I2 => MultOut140, O => Y141, In1IW => Add140aIW, In1FW => Add140aFW, In2IW => Add140bIW, In2FW => Add140bFW);
	WC_Adder141:	WC_AddSub port map (I1 => Y141, I2 => MultOut141, O => Y142, In1IW => Add141aIW, In1FW => Add141aFW, In2IW => Add141bIW, In2FW => Add141bFW);
	WC_Adder142:	WC_AddSub port map (I1 => Y142, I2 => MultOut142, O => Y143, In1IW => Add142aIW, In1FW => Add142aFW, In2IW => Add142bIW, In2FW => Add142bFW);
	WC_Adder143:	WC_AddSub port map (I1 => Y143, I2 => MultOut143, O => Y144, In1IW => Add143aIW, In1FW => Add143aFW, In2IW => Add143bIW, In2FW => Add143bFW);
	WC_Adder144:	WC_AddSub port map (I1 => Y144, I2 => MultOut144, O => Y145, In1IW => Add144aIW, In1FW => Add144aFW, In2IW => Add144bIW, In2FW => Add144bFW);
	WC_Adder145:	WC_AddSub port map (I1 => Y145, I2 => MultOut145, O => Y146, In1IW => Add145aIW, In1FW => Add145aFW, In2IW => Add145bIW, In2FW => Add145bFW);
	WC_Adder146:	WC_AddSub port map (I1 => Y146, I2 => MultOut146, O => Y147, In1IW => Add146aIW, In1FW => Add146aFW, In2IW => Add146bIW, In2FW => Add146bFW);
	WC_Adder147:	WC_AddSub port map (I1 => Y147, I2 => MultOut147, O => Y148, In1IW => Add147aIW, In1FW => Add147aFW, In2IW => Add147bIW, In2FW => Add147bFW);
	WC_Adder148:	WC_AddSub port map (I1 => Y148, I2 => MultOut148, O => Y149, In1IW => Add148aIW, In1FW => Add148aFW, In2IW => Add148bIW, In2FW => Add148bFW);
	WC_Adder149:	WC_AddSub port map (I1 => Y149, I2 => MultOut149, O => Y150, In1IW => Add149aIW, In1FW => Add149aFW, In2IW => Add149bIW, In2FW => Add149bFW);
	WC_Adder150:	WC_AddSub port map (I1 => Y150, I2 => MultOut150, O => Y   , In1IW => Add150aIW, In1FW => Add150aFW, In2IW => Add150bIW, In2FW => Add150bFW);
	

end Behavioral;
